// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : PippengerU250
// Git hash  : fb144932a897c9b17da6701f7d45ebc71bfd9c88

`timescale 1ns/1ps

module PippengerU250 (
  output              dataBus_awvalid,
  input               dataBus_awready,
  output     [63:0]   dataBus_awaddr,
  output     [7:0]    dataBus_awlen,
  output              dataBus_wvalid,
  input               dataBus_wready,
  output     [511:0]  dataBus_wdata,
  output              dataBus_wlast,
  input               dataBus_bvalid,
  output              dataBus_bready,
  output              dataBus_arvalid,
  input               dataBus_arready,
  output     [63:0]   dataBus_araddr,
  output     [7:0]    dataBus_arlen,
  input               dataBus_rvalid,
  output              dataBus_rready,
  input      [511:0]  dataBus_rdata,
  input               dataBus_rlast,
  input               s_axi_control_awvalid,
  output              s_axi_control_awready,
  input      [5:0]    s_axi_control_awaddr,
  input      [2:0]    s_axi_control_awprot,
  input               s_axi_control_wvalid,
  output              s_axi_control_wready,
  input      [31:0]   s_axi_control_wdata,
  input      [3:0]    s_axi_control_wstrb,
  output              s_axi_control_bvalid,
  input               s_axi_control_bready,
  output     [1:0]    s_axi_control_bresp,
  input               s_axi_control_arvalid,
  output reg          s_axi_control_arready,
  input      [5:0]    s_axi_control_araddr,
  input      [2:0]    s_axi_control_arprot,
  output              s_axi_control_rvalid,
  input               s_axi_control_rready,
  output     [31:0]   s_axi_control_rdata,
  output     [1:0]    s_axi_control_rresp,
  input               clk,
  input               resetn
);

  wire       [376:0]  pippenger_1_io_dataIn_payload_fragment_P_X;
  wire       [376:0]  pippenger_1_io_dataIn_payload_fragment_P_Y;
  wire       [376:0]  pippenger_1_io_dataIn_payload_fragment_P_T;
  wire       [252:0]  pippenger_1_io_dataIn_payload_fragment_K;
  wire                dataBusReadArea_inputDMA_io_streamBus_ready;
  wire                pippenger_1_io_dataIn_ready;
  wire                pippenger_1_io_dataOut_valid;
  wire       [376:0]  pippenger_1_io_dataOut_payload_X;
  wire       [376:0]  pippenger_1_io_dataOut_payload_Y;
  wire       [376:0]  pippenger_1_io_dataOut_payload_Z;
  wire       [376:0]  pippenger_1_io_dataOut_payload_T;
  wire                dataBusReadArea_inputDMA_io_axi4Bus_ar_valid;
  wire       [63:0]   dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_addr;
  wire       [7:0]    dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_len;
  wire                dataBusReadArea_inputDMA_io_axi4Bus_r_ready;
  wire                dataBusReadArea_inputDMA_io_streamBus_valid;
  wire       [511:0]  dataBusReadArea_inputDMA_io_streamBus_payload;
  wire                dataBusReadArea_inputDMA_io_done;
  wire       [27:0]   _zz_pageNum;
  wire       [27:0]   _zz_pageNum_1;
  wire       [26:0]   _zz_pageNum_2;
  wire       [26:0]   _zz_pageNum_3;
  wire       [1:0]    _zz_dataBusReadArea_inputCnt_valueNext;
  wire       [0:0]    _zz_dataBusReadArea_inputCnt_valueNext_1;
  wire       [31:0]   _zz_dataBusReadArea_lastCnt_valueNext;
  wire       [0:0]    _zz_dataBusReadArea_lastCnt_valueNext_1;
  wire       [1:0]    _zz_dataBusWriteArea_outputCnt_valueNext;
  wire       [0:0]    _zz_dataBusWriteArea_outputCnt_valueNext_1;
  wire       [376:0]  _zz_dataBus_wdata;
  wire       [31:0]   _zz_startReadAddress;
  wire       [31:0]   _zz_startReadAddress_1;
  wire       [31:0]   _zz_startReadAddress_2;
  wire       [31:0]   _zz_startReadAddress_3;
  wire       [31:0]   _zz_startWriteAddress;
  wire       [31:0]   _zz_startWriteAddress_1;
  wire       [31:0]   _zz_startWriteAddress_2;
  wire       [31:0]   _zz_startWriteAddress_3;
  reg                 startRise;
  reg                 readStart;
  reg                 writeStart;
  reg        [25:0]   num;
  reg        [27:0]   pageNum;
  reg        [63:0]   startReadAddress;
  reg        [63:0]   startWriteAddress;
  wire                slaveFactory_readErrorFlag;
  wire                slaveFactory_writeErrorFlag;
  wire                slaveFactory_readHaltRequest;
  wire                slaveFactory_writeHaltRequest;
  wire                slaveFactory_writeJoinEvent_valid;
  wire                slaveFactory_writeJoinEvent_ready;
  wire                slaveFactory_writeJoinEvent_fire;
  reg        [1:0]    slaveFactory_writeRsp_resp;
  wire                slaveFactory_writeJoinEvent_translated_valid;
  wire                slaveFactory_writeJoinEvent_translated_ready;
  wire       [1:0]    slaveFactory_writeJoinEvent_translated_payload_resp;
  wire                _zz_slaveFactory_writeJoinEvent_translated_ready;
  reg                 _zz_slaveFactory_writeJoinEvent_translated_ready_1;
  wire                _zz_s_axi_control_bvalid;
  reg                 _zz_s_axi_control_bvalid_1;
  reg        [1:0]    _zz_s_axi_control_bresp;
  wire                when_Stream_l368;
  wire                slaveFactory_readDataStage_valid;
  wire                slaveFactory_readDataStage_ready;
  wire       [5:0]    slaveFactory_readDataStage_payload_addr;
  wire       [2:0]    slaveFactory_readDataStage_payload_prot;
  reg                 io_s_axi_control_ar_rValid;
  reg        [5:0]    io_s_axi_control_ar_rData_addr;
  reg        [2:0]    io_s_axi_control_ar_rData_prot;
  wire                when_Stream_l368_1;
  reg        [31:0]   slaveFactory_readRsp_data;
  reg        [1:0]    slaveFactory_readRsp_resp;
  wire                _zz_s_axi_control_rvalid;
  wire       [5:0]    slaveFactory_readAddressMasked;
  wire       [5:0]    slaveFactory_writeAddressMasked;
  wire                slaveFactory_writeOccur;
  wire                slaveFactory_readOccur;
  wire       [63:0]   _zz_slaveFactory_readRsp_data;
  wire       [63:0]   _zz_slaveFactory_readRsp_data_1;
  reg                 dataBusReadArea_inputCnt_willIncrement;
  wire                dataBusReadArea_inputCnt_willClear;
  reg        [1:0]    dataBusReadArea_inputCnt_valueNext;
  reg        [1:0]    dataBusReadArea_inputCnt_value;
  reg                 dataBusReadArea_inputCnt_willOverflowIfInc;
  wire                dataBusReadArea_inputCnt_willOverflow;
  reg                 dataBusReadArea_inputValid;
  reg        [511:0]  dataBusReadArea_inputData_0;
  reg        [511:0]  dataBusReadArea_inputData_1;
  reg        [511:0]  dataBusReadArea_inputData_2;
  wire       [383:0]  dataBusReadArea_outputData_0;
  wire       [383:0]  dataBusReadArea_outputData_1;
  wire       [383:0]  dataBusReadArea_outputData_2;
  wire       [383:0]  dataBusReadArea_outputData_3;
  wire       [1535:0] _zz_dataBusReadArea_outputData_0;
  reg                 dataBusReadArea_lastCnt_willIncrement;
  reg                 dataBusReadArea_lastCnt_willClear;
  reg        [31:0]   dataBusReadArea_lastCnt_valueNext;
  reg        [31:0]   dataBusReadArea_lastCnt_value;
  reg                 dataBusReadArea_lastCnt_willOverflowIfInc;
  wire                dataBusReadArea_lastCnt_willOverflow;
  wire                toplevel_pippenger_1_io_dataIn_fire;
  reg                 _zz_1;
  reg                 _zz_io_dataIn_payload_last;
  wire                toplevel_dataBusReadArea_inputDMA_io_streamBus_fire;
  reg                 dataBusWriteArea_outputCnt_willIncrement;
  wire                dataBusWriteArea_outputCnt_willClear;
  reg        [1:0]    dataBusWriteArea_outputCnt_valueNext;
  reg        [1:0]    dataBusWriteArea_outputCnt_value;
  reg                 dataBusWriteArea_outputCnt_willOverflowIfInc;
  wire                dataBusWriteArea_outputCnt_willOverflow;
  reg                 dataBusWriteArea_dataOutputValid;
  reg        [376:0]  dataBusWriteArea_dataReg_0;
  reg        [376:0]  dataBusWriteArea_dataReg_1;
  reg        [376:0]  dataBusWriteArea_dataReg_2;
  reg        [376:0]  dataBusWriteArea_dataReg_3;
  reg                 dataBusWriteArea_addressOutputValid;
  wire                io_dataBus_w_fire;
  wire                when_AxiLite4SlaveFactory_l68;
  wire                when_AxiLite4SlaveFactory_l68_1;
  wire                when_AxiLite4SlaveFactory_l68_2;
  wire                when_AxiLite4SlaveFactory_l68_3;
  wire                when_AxiLite4SlaveFactory_l86;
  wire                when_AxiLite4SlaveFactory_l86_1;
  wire                when_AxiLite4SlaveFactory_l86_2;
  wire                when_AxiLite4SlaveFactory_l86_3;

  assign _zz_pageNum = (_zz_pageNum_1 + {1'b0,_zz_pageNum_3});
  assign _zz_pageNum_2 = {1'b0,num};
  assign _zz_pageNum_1 = {1'd0, _zz_pageNum_2};
  assign _zz_pageNum_3 = ({1'd0,num} <<< 1);
  assign _zz_dataBusReadArea_inputCnt_valueNext_1 = dataBusReadArea_inputCnt_willIncrement;
  assign _zz_dataBusReadArea_inputCnt_valueNext = {1'd0, _zz_dataBusReadArea_inputCnt_valueNext_1};
  assign _zz_dataBusReadArea_lastCnt_valueNext_1 = dataBusReadArea_lastCnt_willIncrement;
  assign _zz_dataBusReadArea_lastCnt_valueNext = {31'd0, _zz_dataBusReadArea_lastCnt_valueNext_1};
  assign _zz_dataBusWriteArea_outputCnt_valueNext_1 = dataBusWriteArea_outputCnt_willIncrement;
  assign _zz_dataBusWriteArea_outputCnt_valueNext = {1'd0, _zz_dataBusWriteArea_outputCnt_valueNext_1};
  assign _zz_dataBus_wdata = dataBusWriteArea_dataReg_0;
  assign _zz_startReadAddress_1 = s_axi_control_wdata[31 : 0];
  assign _zz_startReadAddress = _zz_startReadAddress_1;
  assign _zz_startReadAddress_3 = s_axi_control_wdata[31 : 0];
  assign _zz_startReadAddress_2 = _zz_startReadAddress_3;
  assign _zz_startWriteAddress_1 = s_axi_control_wdata[31 : 0];
  assign _zz_startWriteAddress = _zz_startWriteAddress_1;
  assign _zz_startWriteAddress_3 = s_axi_control_wdata[31 : 0];
  assign _zz_startWriteAddress_2 = _zz_startWriteAddress_3;
  PippengerWithPAdd pippenger_1 (
    .io_dataIn_valid                (dataBusReadArea_inputValid                                                                          ), //i
    .io_dataIn_ready                (pippenger_1_io_dataIn_ready                                                                         ), //o
    .io_dataIn_payload_last         (_zz_io_dataIn_payload_last                                                                          ), //i
    .io_dataIn_payload_fragment_P_X (pippenger_1_io_dataIn_payload_fragment_P_X[376:0]                                                   ), //i
    .io_dataIn_payload_fragment_P_Y (pippenger_1_io_dataIn_payload_fragment_P_Y[376:0]                                                   ), //i
    .io_dataIn_payload_fragment_P_Z (377'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001), //i
    .io_dataIn_payload_fragment_P_T (pippenger_1_io_dataIn_payload_fragment_P_T[376:0]                                                   ), //i
    .io_dataIn_payload_fragment_K   (pippenger_1_io_dataIn_payload_fragment_K[252:0]                                                     ), //i
    .io_dataOut_valid               (pippenger_1_io_dataOut_valid                                                                        ), //o
    .io_dataOut_ready               (1'b1                                                                                                ), //i
    .io_dataOut_payload_X           (pippenger_1_io_dataOut_payload_X[376:0]                                                             ), //o
    .io_dataOut_payload_Y           (pippenger_1_io_dataOut_payload_Y[376:0]                                                             ), //o
    .io_dataOut_payload_Z           (pippenger_1_io_dataOut_payload_Z[376:0]                                                             ), //o
    .io_dataOut_payload_T           (pippenger_1_io_dataOut_payload_T[376:0]                                                             ), //o
    .clk                            (clk                                                                                                 ), //i
    .resetn                         (resetn                                                                                              )  //i
  );
  Axi4PageRDMA dataBusReadArea_inputDMA (
    .io_axi4Bus_ar_valid        (dataBusReadArea_inputDMA_io_axi4Bus_ar_valid             ), //o
    .io_axi4Bus_ar_ready        (dataBus_arready                                          ), //i
    .io_axi4Bus_ar_payload_addr (dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_addr[63:0]), //o
    .io_axi4Bus_ar_payload_len  (dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_len[7:0]  ), //o
    .io_axi4Bus_r_valid         (dataBus_rvalid                                           ), //i
    .io_axi4Bus_r_ready         (dataBusReadArea_inputDMA_io_axi4Bus_r_ready              ), //o
    .io_axi4Bus_r_payload_data  (dataBus_rdata[511:0]                                     ), //i
    .io_axi4Bus_r_payload_last  (dataBus_rlast                                            ), //i
    .io_streamBus_valid         (dataBusReadArea_inputDMA_io_streamBus_valid              ), //o
    .io_streamBus_ready         (dataBusReadArea_inputDMA_io_streamBus_ready              ), //i
    .io_streamBus_payload       (dataBusReadArea_inputDMA_io_streamBus_payload[511:0]     ), //o
    .io_work                    (readStart                                                ), //i
    .io_address                 (startReadAddress[63:0]                                   ), //i
    .io_pageNum                 (pageNum[27:0]                                            ), //i
    .io_done                    (dataBusReadArea_inputDMA_io_done                         ), //o
    .clk                        (clk                                                      ), //i
    .resetn                     (resetn                                                   )  //i
  );
  always @(*) begin
    startRise = 1'b0;
    case(slaveFactory_writeAddressMasked)
      6'h10 : begin
        if(slaveFactory_writeOccur) begin
          startRise = s_axi_control_wdata[0];
        end
      end
      default : begin
      end
    endcase
  end

  assign slaveFactory_readErrorFlag = 1'b0;
  assign slaveFactory_writeErrorFlag = 1'b0;
  assign slaveFactory_readHaltRequest = 1'b0;
  assign slaveFactory_writeHaltRequest = 1'b0;
  assign slaveFactory_writeJoinEvent_fire = (slaveFactory_writeJoinEvent_valid && slaveFactory_writeJoinEvent_ready);
  assign slaveFactory_writeJoinEvent_valid = (s_axi_control_awvalid && s_axi_control_wvalid);
  assign s_axi_control_awready = slaveFactory_writeJoinEvent_fire;
  assign s_axi_control_wready = slaveFactory_writeJoinEvent_fire;
  assign slaveFactory_writeJoinEvent_translated_valid = slaveFactory_writeJoinEvent_valid;
  assign slaveFactory_writeJoinEvent_ready = slaveFactory_writeJoinEvent_translated_ready;
  assign slaveFactory_writeJoinEvent_translated_payload_resp = slaveFactory_writeRsp_resp;
  assign _zz_slaveFactory_writeJoinEvent_translated_ready = (! slaveFactory_writeHaltRequest);
  assign slaveFactory_writeJoinEvent_translated_ready = (_zz_slaveFactory_writeJoinEvent_translated_ready_1 && _zz_slaveFactory_writeJoinEvent_translated_ready);
  always @(*) begin
    _zz_slaveFactory_writeJoinEvent_translated_ready_1 = s_axi_control_bready;
    if(when_Stream_l368) begin
      _zz_slaveFactory_writeJoinEvent_translated_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l368 = (! _zz_s_axi_control_bvalid);
  assign _zz_s_axi_control_bvalid = _zz_s_axi_control_bvalid_1;
  assign s_axi_control_bvalid = _zz_s_axi_control_bvalid;
  assign s_axi_control_bresp = _zz_s_axi_control_bresp;
  always @(*) begin
    s_axi_control_arready = slaveFactory_readDataStage_ready;
    if(when_Stream_l368_1) begin
      s_axi_control_arready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! slaveFactory_readDataStage_valid);
  assign slaveFactory_readDataStage_valid = io_s_axi_control_ar_rValid;
  assign slaveFactory_readDataStage_payload_addr = io_s_axi_control_ar_rData_addr;
  assign slaveFactory_readDataStage_payload_prot = io_s_axi_control_ar_rData_prot;
  assign _zz_s_axi_control_rvalid = (! slaveFactory_readHaltRequest);
  assign slaveFactory_readDataStage_ready = (s_axi_control_rready && _zz_s_axi_control_rvalid);
  assign s_axi_control_rvalid = (slaveFactory_readDataStage_valid && _zz_s_axi_control_rvalid);
  assign s_axi_control_rdata = slaveFactory_readRsp_data;
  assign s_axi_control_rresp = slaveFactory_readRsp_resp;
  always @(*) begin
    if(slaveFactory_writeErrorFlag) begin
      slaveFactory_writeRsp_resp = 2'b10;
    end else begin
      slaveFactory_writeRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    if(slaveFactory_readErrorFlag) begin
      slaveFactory_readRsp_resp = 2'b10;
    end else begin
      slaveFactory_readRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    slaveFactory_readRsp_data = 32'h0;
    case(slaveFactory_readAddressMasked)
      6'h10 : begin
        slaveFactory_readRsp_data[0 : 0] = (readStart || writeStart);
      end
      6'h18 : begin
        slaveFactory_readRsp_data[31 : 0] = {num,6'h3f};
      end
      default : begin
      end
    endcase
    if(when_AxiLite4SlaveFactory_l86) begin
      slaveFactory_readRsp_data[31 : 0] = _zz_slaveFactory_readRsp_data[31 : 0];
    end
    if(when_AxiLite4SlaveFactory_l86_1) begin
      slaveFactory_readRsp_data[31 : 0] = _zz_slaveFactory_readRsp_data[63 : 32];
    end
    if(when_AxiLite4SlaveFactory_l86_2) begin
      slaveFactory_readRsp_data[31 : 0] = _zz_slaveFactory_readRsp_data_1[31 : 0];
    end
    if(when_AxiLite4SlaveFactory_l86_3) begin
      slaveFactory_readRsp_data[31 : 0] = _zz_slaveFactory_readRsp_data_1[63 : 32];
    end
  end

  assign slaveFactory_readAddressMasked = (slaveFactory_readDataStage_payload_addr & (~ 6'h03));
  assign slaveFactory_writeAddressMasked = (s_axi_control_awaddr & (~ 6'h03));
  assign slaveFactory_writeOccur = (slaveFactory_writeJoinEvent_valid && slaveFactory_writeJoinEvent_ready);
  assign slaveFactory_readOccur = (s_axi_control_rvalid && s_axi_control_rready);
  assign _zz_slaveFactory_readRsp_data = startReadAddress;
  assign _zz_slaveFactory_readRsp_data_1 = startWriteAddress;
  assign dataBus_arvalid = dataBusReadArea_inputDMA_io_axi4Bus_ar_valid;
  assign dataBus_araddr = dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_addr;
  assign dataBus_arlen = dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_len;
  assign dataBus_rready = dataBusReadArea_inputDMA_io_axi4Bus_r_ready;
  always @(*) begin
    dataBusReadArea_inputCnt_willIncrement = 1'b0;
    if(toplevel_dataBusReadArea_inputDMA_io_streamBus_fire) begin
      dataBusReadArea_inputCnt_willIncrement = 1'b1;
    end
  end

  assign dataBusReadArea_inputCnt_willClear = 1'b0;
  assign dataBusReadArea_inputCnt_willOverflow = (dataBusReadArea_inputCnt_willOverflowIfInc && dataBusReadArea_inputCnt_willIncrement);
  always @(*) begin
    if(dataBusReadArea_inputCnt_willOverflow) begin
      dataBusReadArea_inputCnt_valueNext = 2'b00;
    end else begin
      dataBusReadArea_inputCnt_valueNext = (dataBusReadArea_inputCnt_value + _zz_dataBusReadArea_inputCnt_valueNext);
    end
    if(dataBusReadArea_inputCnt_willClear) begin
      dataBusReadArea_inputCnt_valueNext = 2'b00;
    end
  end

  assign _zz_dataBusReadArea_outputData_0 = {dataBusReadArea_inputData_2,{dataBusReadArea_inputData_1,dataBusReadArea_inputData_0}};
  assign dataBusReadArea_outputData_0 = _zz_dataBusReadArea_outputData_0[383 : 0];
  assign dataBusReadArea_outputData_1 = _zz_dataBusReadArea_outputData_0[767 : 384];
  assign dataBusReadArea_outputData_2 = _zz_dataBusReadArea_outputData_0[1151 : 768];
  assign dataBusReadArea_outputData_3 = _zz_dataBusReadArea_outputData_0[1535 : 1152];
  always @(*) begin
    dataBusReadArea_lastCnt_willIncrement = 1'b0;
    if(toplevel_pippenger_1_io_dataIn_fire) begin
      dataBusReadArea_lastCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    dataBusReadArea_lastCnt_willClear = 1'b0;
    if(toplevel_pippenger_1_io_dataIn_fire) begin
      if(_zz_1) begin
        dataBusReadArea_lastCnt_willClear = 1'b1;
      end
    end
  end

  assign dataBusReadArea_lastCnt_willOverflow = (dataBusReadArea_lastCnt_willOverflowIfInc && dataBusReadArea_lastCnt_willIncrement);
  always @(*) begin
    dataBusReadArea_lastCnt_valueNext = (dataBusReadArea_lastCnt_value + _zz_dataBusReadArea_lastCnt_valueNext);
    if(dataBusReadArea_lastCnt_willClear) begin
      dataBusReadArea_lastCnt_valueNext = 32'h0;
    end
  end

  assign toplevel_pippenger_1_io_dataIn_fire = (dataBusReadArea_inputValid && pippenger_1_io_dataIn_ready);
  assign pippenger_1_io_dataIn_payload_fragment_P_X = dataBusReadArea_outputData_0[376:0];
  assign pippenger_1_io_dataIn_payload_fragment_P_Y = dataBusReadArea_outputData_1[376:0];
  assign pippenger_1_io_dataIn_payload_fragment_P_T = dataBusReadArea_outputData_2[376:0];
  assign pippenger_1_io_dataIn_payload_fragment_K = dataBusReadArea_outputData_3[252:0];
  assign dataBusReadArea_inputDMA_io_streamBus_ready = ((! dataBusReadArea_inputValid) || pippenger_1_io_dataIn_ready);
  assign toplevel_dataBusReadArea_inputDMA_io_streamBus_fire = (dataBusReadArea_inputDMA_io_streamBus_valid && dataBusReadArea_inputDMA_io_streamBus_ready);
  always @(*) begin
    dataBusWriteArea_outputCnt_willIncrement = 1'b0;
    if(io_dataBus_w_fire) begin
      dataBusWriteArea_outputCnt_willIncrement = 1'b1;
    end
  end

  assign dataBusWriteArea_outputCnt_willClear = 1'b0;
  assign dataBusWriteArea_outputCnt_willOverflow = (dataBusWriteArea_outputCnt_willOverflowIfInc && dataBusWriteArea_outputCnt_willIncrement);
  always @(*) begin
    dataBusWriteArea_outputCnt_valueNext = (dataBusWriteArea_outputCnt_value + _zz_dataBusWriteArea_outputCnt_valueNext);
    if(dataBusWriteArea_outputCnt_willClear) begin
      dataBusWriteArea_outputCnt_valueNext = 2'b00;
    end
  end

  assign dataBus_awvalid = dataBusWriteArea_addressOutputValid;
  assign dataBus_awaddr = startWriteAddress;
  assign dataBus_awlen = 8'h03;
  assign dataBus_wvalid = dataBusWriteArea_dataOutputValid;
  assign dataBus_wdata = {135'd0, _zz_dataBus_wdata};
  assign dataBus_wlast = dataBusWriteArea_outputCnt_willOverflowIfInc;
  assign io_dataBus_w_fire = (dataBus_wvalid && dataBus_wready);
  assign dataBus_bready = 1'b1;
  assign when_AxiLite4SlaveFactory_l68 = ((slaveFactory_writeAddressMasked & (~ 6'h03)) == 6'h20);
  assign when_AxiLite4SlaveFactory_l68_1 = ((slaveFactory_writeAddressMasked & (~ 6'h03)) == 6'h24);
  assign when_AxiLite4SlaveFactory_l68_2 = ((slaveFactory_writeAddressMasked & (~ 6'h03)) == 6'h28);
  assign when_AxiLite4SlaveFactory_l68_3 = ((slaveFactory_writeAddressMasked & (~ 6'h03)) == 6'h2c);
  assign when_AxiLite4SlaveFactory_l86 = ((slaveFactory_readAddressMasked & (~ 6'h03)) == 6'h20);
  assign when_AxiLite4SlaveFactory_l86_1 = ((slaveFactory_readAddressMasked & (~ 6'h03)) == 6'h24);
  assign when_AxiLite4SlaveFactory_l86_2 = ((slaveFactory_readAddressMasked & (~ 6'h03)) == 6'h28);
  assign when_AxiLite4SlaveFactory_l86_3 = ((slaveFactory_readAddressMasked & (~ 6'h03)) == 6'h2c);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      readStart <= 1'b0;
      writeStart <= 1'b0;
      _zz_s_axi_control_bvalid_1 <= 1'b0;
      io_s_axi_control_ar_rValid <= 1'b0;
      dataBusReadArea_inputCnt_value <= 2'b00;
      dataBusReadArea_inputCnt_willOverflowIfInc <= 1'b0;
      dataBusReadArea_inputValid <= 1'b0;
      dataBusReadArea_lastCnt_value <= 32'h0;
      dataBusReadArea_lastCnt_willOverflowIfInc <= 1'b0;
      dataBusWriteArea_outputCnt_value <= 2'b00;
      dataBusWriteArea_outputCnt_willOverflowIfInc <= 1'b0;
      dataBusWriteArea_dataOutputValid <= 1'b0;
      dataBusWriteArea_addressOutputValid <= 1'b0;
    end else begin
      if(startRise) begin
        readStart <= 1'b1;
      end
      if(startRise) begin
        writeStart <= 1'b1;
      end
      if(_zz_slaveFactory_writeJoinEvent_translated_ready_1) begin
        _zz_s_axi_control_bvalid_1 <= (slaveFactory_writeJoinEvent_translated_valid && _zz_slaveFactory_writeJoinEvent_translated_ready);
      end
      if(s_axi_control_arready) begin
        io_s_axi_control_ar_rValid <= s_axi_control_arvalid;
      end
      if(dataBusReadArea_inputDMA_io_done) begin
        readStart <= 1'b0;
      end
      dataBusReadArea_inputCnt_value <= dataBusReadArea_inputCnt_valueNext;
      dataBusReadArea_inputCnt_willOverflowIfInc <= (dataBusReadArea_inputCnt_valueNext == 2'b10);
      dataBusReadArea_lastCnt_value <= dataBusReadArea_lastCnt_valueNext;
      dataBusReadArea_lastCnt_willOverflowIfInc <= (dataBusReadArea_lastCnt_valueNext == 32'hffffffff);
      if(dataBusReadArea_inputCnt_willOverflow) begin
        dataBusReadArea_inputValid <= 1'b1;
      end else begin
        if(pippenger_1_io_dataIn_ready) begin
          dataBusReadArea_inputValid <= 1'b0;
        end
      end
      dataBusWriteArea_outputCnt_value <= dataBusWriteArea_outputCnt_valueNext;
      dataBusWriteArea_outputCnt_willOverflowIfInc <= (dataBusWriteArea_outputCnt_valueNext == 2'b11);
      if(pippenger_1_io_dataOut_valid) begin
        dataBusWriteArea_dataOutputValid <= 1'b1;
      end else begin
        if(dataBusWriteArea_outputCnt_willOverflow) begin
          dataBusWriteArea_dataOutputValid <= 1'b0;
        end
      end
      if(pippenger_1_io_dataOut_valid) begin
        dataBusWriteArea_addressOutputValid <= 1'b1;
      end else begin
        if(dataBus_arready) begin
          dataBusWriteArea_addressOutputValid <= 1'b0;
        end
      end
      if(dataBus_bvalid) begin
        writeStart <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    pageNum <= (_zz_pageNum + 28'h0000002);
    if(_zz_slaveFactory_writeJoinEvent_translated_ready_1) begin
      _zz_s_axi_control_bresp <= slaveFactory_writeJoinEvent_translated_payload_resp;
    end
    if(s_axi_control_arready) begin
      io_s_axi_control_ar_rData_addr <= s_axi_control_araddr;
      io_s_axi_control_ar_rData_prot <= s_axi_control_arprot;
    end
    _zz_io_dataIn_payload_last <= (dataBusReadArea_lastCnt_valueNext == {num,6'h3f});
    if(toplevel_dataBusReadArea_inputDMA_io_streamBus_fire) begin
      dataBusReadArea_inputData_0 <= dataBusReadArea_inputData_1;
      dataBusReadArea_inputData_1 <= dataBusReadArea_inputData_2;
      dataBusReadArea_inputData_2 <= dataBusReadArea_inputDMA_io_streamBus_payload;
    end
    if(pippenger_1_io_dataOut_valid) begin
      dataBusWriteArea_dataReg_0 <= pippenger_1_io_dataOut_payload_X;
      dataBusWriteArea_dataReg_1 <= pippenger_1_io_dataOut_payload_Y;
      dataBusWriteArea_dataReg_2 <= pippenger_1_io_dataOut_payload_Z;
      dataBusWriteArea_dataReg_3 <= pippenger_1_io_dataOut_payload_T;
    end else begin
      if(dataBus_wready) begin
        dataBusWriteArea_dataReg_0 <= dataBusWriteArea_dataReg_1;
        dataBusWriteArea_dataReg_1 <= dataBusWriteArea_dataReg_2;
        dataBusWriteArea_dataReg_2 <= dataBusWriteArea_dataReg_3;
      end
    end
    case(slaveFactory_writeAddressMasked)
      6'h18 : begin
        if(slaveFactory_writeOccur) begin
          num <= s_axi_control_wdata[31 : 6];
        end
      end
      default : begin
      end
    endcase
    if(when_AxiLite4SlaveFactory_l68) begin
      if(slaveFactory_writeOccur) begin
        startReadAddress[31 : 0] <= _zz_startReadAddress;
      end
    end
    if(when_AxiLite4SlaveFactory_l68_1) begin
      if(slaveFactory_writeOccur) begin
        startReadAddress[63 : 32] <= _zz_startReadAddress_2;
      end
    end
    if(when_AxiLite4SlaveFactory_l68_2) begin
      if(slaveFactory_writeOccur) begin
        startWriteAddress[31 : 0] <= _zz_startWriteAddress;
      end
    end
    if(when_AxiLite4SlaveFactory_l68_3) begin
      if(slaveFactory_writeOccur) begin
        startWriteAddress[63 : 32] <= _zz_startWriteAddress_2;
      end
    end
  end

  always @(posedge clk) begin
    _zz_1 <= (dataBusReadArea_lastCnt_valueNext == {num,6'h3f});
  end


endmodule

module Axi4PageRDMA (
  output reg          io_axi4Bus_ar_valid,
  input               io_axi4Bus_ar_ready,
  output reg [63:0]   io_axi4Bus_ar_payload_addr,
  output reg [7:0]    io_axi4Bus_ar_payload_len,
  input               io_axi4Bus_r_valid,
  output              io_axi4Bus_r_ready,
  input      [511:0]  io_axi4Bus_r_payload_data,
  input               io_axi4Bus_r_payload_last,
  output              io_streamBus_valid,
  input               io_streamBus_ready,
  output     [511:0]  io_streamBus_payload,
  input               io_work,
  input      [63:0]   io_address,
  input      [27:0]   io_pageNum,
  output reg          io_done,
  input               clk,
  input               resetn
);

  wire                readFifo_io_push_ready;
  wire                readFifo_io_pop_valid;
  wire       [511:0]  readFifo_io_pop_payload;
  wire       [7:0]    readFifo_io_pushPtr;
  wire       [7:0]    readFifo_io_popPtr;
  wire       [27:0]   _zz_readArea_addressCnt_valueNext;
  wire       [0:0]    _zz_readArea_addressCnt_valueNext_1;
  wire       [1:0]    _zz_readArea_outStandingCnt_valueNext;
  wire       [0:0]    _zz_readArea_outStandingCnt_valueNext_1;
  wire       [51:0]   _zz_io_axi4Bus_ar_payload_addr;
  wire       [51:0]   _zz_io_axi4Bus_ar_payload_addr_1;
  wire                io_axi4Bus_r_translated_valid;
  wire                io_axi4Bus_r_translated_ready;
  wire       [511:0]  io_axi4Bus_r_translated_payload;
  reg                 readArea_addressCnt_willIncrement;
  reg                 readArea_addressCnt_willClear;
  reg        [27:0]   readArea_addressCnt_valueNext;
  reg        [27:0]   readArea_addressCnt_value;
  reg                 readArea_addressCnt_willOverflowIfInc;
  wire                readArea_addressCnt_willOverflow;
  reg                 readArea_outStandingCnt_willIncrement;
  wire                readArea_outStandingCnt_willClear;
  reg        [1:0]    readArea_outStandingCnt_valueNext;
  reg        [1:0]    readArea_outStandingCnt_value;
  reg                 readArea_outStandingCnt_willOverflowIfInc;
  wire                readArea_outStandingCnt_willOverflow;
  wire       [1:0]    _zz_io_axi4Bus_ar_valid;
  reg                 _zz_io_axi4Bus_ar_valid_1;
  wire                io_axi4Bus_ar_fire;
  reg                 _zz_1;

  assign _zz_readArea_addressCnt_valueNext_1 = readArea_addressCnt_willIncrement;
  assign _zz_readArea_addressCnt_valueNext = {27'd0, _zz_readArea_addressCnt_valueNext_1};
  assign _zz_readArea_outStandingCnt_valueNext_1 = readArea_outStandingCnt_willIncrement;
  assign _zz_readArea_outStandingCnt_valueNext = {1'd0, _zz_readArea_outStandingCnt_valueNext_1};
  assign _zz_io_axi4Bus_ar_payload_addr = (io_address[63 : 12] + _zz_io_axi4Bus_ar_payload_addr_1);
  assign _zz_io_axi4Bus_ar_payload_addr_1 = {24'd0, readArea_addressCnt_value};
  FIFO readFifo (
    .io_push_valid   (io_axi4Bus_r_translated_valid         ), //i
    .io_push_ready   (readFifo_io_push_ready                ), //o
    .io_push_payload (io_axi4Bus_r_translated_payload[511:0]), //i
    .io_pop_valid    (readFifo_io_pop_valid                 ), //o
    .io_pop_ready    (io_streamBus_ready                    ), //i
    .io_pop_payload  (readFifo_io_pop_payload[511:0]        ), //o
    .io_pushPtr      (readFifo_io_pushPtr[7:0]              ), //o
    .io_popPtr       (readFifo_io_popPtr[7:0]               ), //o
    .clk             (clk                                   ), //i
    .resetn          (resetn                                )  //i
  );
  assign io_streamBus_valid = readFifo_io_pop_valid;
  assign io_streamBus_payload = readFifo_io_pop_payload;
  assign io_axi4Bus_r_translated_valid = io_axi4Bus_r_valid;
  assign io_axi4Bus_r_ready = io_axi4Bus_r_translated_ready;
  assign io_axi4Bus_r_translated_payload = io_axi4Bus_r_payload_data;
  assign io_axi4Bus_r_translated_ready = readFifo_io_push_ready;
  always @(*) begin
    readArea_addressCnt_willIncrement = 1'b0;
    if(io_axi4Bus_ar_fire) begin
      readArea_addressCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    readArea_addressCnt_willClear = 1'b0;
    if(io_axi4Bus_ar_fire) begin
      if(_zz_1) begin
        readArea_addressCnt_willClear = 1'b1;
      end
    end
  end

  assign readArea_addressCnt_willOverflow = (readArea_addressCnt_willOverflowIfInc && readArea_addressCnt_willIncrement);
  always @(*) begin
    readArea_addressCnt_valueNext = (readArea_addressCnt_value + _zz_readArea_addressCnt_valueNext);
    if(readArea_addressCnt_willClear) begin
      readArea_addressCnt_valueNext = 28'h0;
    end
  end

  always @(*) begin
    readArea_outStandingCnt_willIncrement = 1'b0;
    if(io_axi4Bus_ar_fire) begin
      readArea_outStandingCnt_willIncrement = 1'b1;
    end
  end

  assign readArea_outStandingCnt_willClear = 1'b0;
  assign readArea_outStandingCnt_willOverflow = (readArea_outStandingCnt_willOverflowIfInc && readArea_outStandingCnt_willIncrement);
  always @(*) begin
    readArea_outStandingCnt_valueNext = (readArea_outStandingCnt_value + _zz_readArea_outStandingCnt_valueNext);
    if(readArea_outStandingCnt_willClear) begin
      readArea_outStandingCnt_valueNext = 2'b00;
    end
  end

  always @(*) begin
    io_axi4Bus_ar_valid = 1'b0;
    if(io_work) begin
      io_axi4Bus_ar_valid = _zz_io_axi4Bus_ar_valid_1;
    end
  end

  always @(*) begin
    io_axi4Bus_ar_payload_addr = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(io_work) begin
      io_axi4Bus_ar_payload_addr = {_zz_io_axi4Bus_ar_payload_addr,12'h0};
    end
  end

  always @(*) begin
    io_axi4Bus_ar_payload_len = 8'bxxxxxxxx;
    if(io_work) begin
      io_axi4Bus_ar_payload_len = 8'h3f;
    end
  end

  always @(*) begin
    io_done = 1'b0;
    if(io_axi4Bus_ar_fire) begin
      if(_zz_1) begin
        io_done = 1'b1;
      end
    end
  end

  assign _zz_io_axi4Bus_ar_valid = readFifo_io_popPtr[7 : 6];
  assign io_axi4Bus_ar_fire = (io_axi4Bus_ar_valid && io_axi4Bus_ar_ready);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      readArea_addressCnt_value <= 28'h0;
      readArea_addressCnt_willOverflowIfInc <= 1'b0;
      readArea_outStandingCnt_value <= 2'b00;
      readArea_outStandingCnt_willOverflowIfInc <= 1'b0;
    end else begin
      readArea_addressCnt_value <= readArea_addressCnt_valueNext;
      readArea_addressCnt_willOverflowIfInc <= (readArea_addressCnt_valueNext == 28'hfffffff);
      readArea_outStandingCnt_value <= readArea_outStandingCnt_valueNext;
      readArea_outStandingCnt_willOverflowIfInc <= (readArea_outStandingCnt_valueNext == 2'b11);
    end
  end

  always @(posedge clk) begin
    _zz_io_axi4Bus_ar_valid_1 <= (! ((readArea_outStandingCnt_valueNext[1] != _zz_io_axi4Bus_ar_valid[1]) && (readArea_outStandingCnt_valueNext[0 : 0] == _zz_io_axi4Bus_ar_valid[0 : 0])));
  end

  always @(posedge clk) begin
    _zz_1 <= (readArea_addressCnt_valueNext == io_pageNum);
  end


endmodule

module PippengerWithPAdd (
  input               io_dataIn_valid,
  output              io_dataIn_ready,
  input               io_dataIn_payload_last,
  input      [376:0]  io_dataIn_payload_fragment_P_X,
  input      [376:0]  io_dataIn_payload_fragment_P_Y,
  input      [376:0]  io_dataIn_payload_fragment_P_Z,
  input      [376:0]  io_dataIn_payload_fragment_P_T,
  input      [252:0]  io_dataIn_payload_fragment_K,
  output              io_dataOut_valid,
  input               io_dataOut_ready,
  output     [376:0]  io_dataOut_payload_X,
  output     [376:0]  io_dataOut_payload_Y,
  output     [376:0]  io_dataOut_payload_Z,
  output     [376:0]  io_dataOut_payload_T,
  input               clk,
  input               resetn
);

  wire       [376:0]  adder_0_io_s_X;
  wire       [376:0]  adder_0_io_s_Y;
  wire       [376:0]  adder_0_io_s_Z;
  wire       [376:0]  adder_0_io_s_T;
  wire       [376:0]  adder_1_io_s_X;
  wire       [376:0]  adder_1_io_s_Y;
  wire       [376:0]  adder_1_io_s_Z;
  wire       [376:0]  adder_1_io_s_T;
  wire       [376:0]  neg_io_n_X;
  wire       [376:0]  neg_io_n_Y;
  wire       [376:0]  neg_io_n_Z;
  wire       [376:0]  neg_io_n_T;
  wire                pippenger_1_io_dataIn_ready;
  wire                pippenger_1_io_dataOut_valid;
  wire       [376:0]  pippenger_1_io_dataOut_payload_X;
  wire       [376:0]  pippenger_1_io_dataOut_payload_Y;
  wire       [376:0]  pippenger_1_io_dataOut_payload_Z;
  wire       [376:0]  pippenger_1_io_dataOut_payload_T;
  wire       [376:0]  pippenger_1_pAddPort_0_a_X;
  wire       [376:0]  pippenger_1_pAddPort_0_a_Y;
  wire       [376:0]  pippenger_1_pAddPort_0_a_Z;
  wire       [376:0]  pippenger_1_pAddPort_0_a_T;
  wire       [376:0]  pippenger_1_pAddPort_0_b_X;
  wire       [376:0]  pippenger_1_pAddPort_0_b_Y;
  wire       [376:0]  pippenger_1_pAddPort_0_b_Z;
  wire       [376:0]  pippenger_1_pAddPort_0_b_T;
  wire       [376:0]  pippenger_1_pAddPort_1_a_X;
  wire       [376:0]  pippenger_1_pAddPort_1_a_Y;
  wire       [376:0]  pippenger_1_pAddPort_1_a_Z;
  wire       [376:0]  pippenger_1_pAddPort_1_a_T;
  wire       [376:0]  pippenger_1_pAddPort_1_b_X;
  wire       [376:0]  pippenger_1_pAddPort_1_b_Y;
  wire       [376:0]  pippenger_1_pAddPort_1_b_Z;
  wire       [376:0]  pippenger_1_pAddPort_1_b_T;
  wire       [376:0]  pippenger_1_pNegPort_a_X;
  wire       [376:0]  pippenger_1_pNegPort_a_Y;
  wire       [376:0]  pippenger_1_pNegPort_a_Z;
  wire       [376:0]  pippenger_1_pNegPort_a_T;

  PAdd adder_0 (
    .io_a_X (pippenger_1_pAddPort_0_a_X[376:0]), //i
    .io_a_Y (pippenger_1_pAddPort_0_a_Y[376:0]), //i
    .io_a_Z (pippenger_1_pAddPort_0_a_Z[376:0]), //i
    .io_a_T (pippenger_1_pAddPort_0_a_T[376:0]), //i
    .io_b_X (pippenger_1_pAddPort_0_b_X[376:0]), //i
    .io_b_Y (pippenger_1_pAddPort_0_b_Y[376:0]), //i
    .io_b_Z (pippenger_1_pAddPort_0_b_Z[376:0]), //i
    .io_b_T (pippenger_1_pAddPort_0_b_T[376:0]), //i
    .io_s_X (adder_0_io_s_X[376:0]            ), //o
    .io_s_Y (adder_0_io_s_Y[376:0]            ), //o
    .io_s_Z (adder_0_io_s_Z[376:0]            ), //o
    .io_s_T (adder_0_io_s_T[376:0]            ), //o
    .clk    (clk                              ), //i
    .resetn (resetn                           )  //i
  );
  PAdd_1 adder_1 (
    .io_a_X (pippenger_1_pAddPort_1_a_X[376:0]), //i
    .io_a_Y (pippenger_1_pAddPort_1_a_Y[376:0]), //i
    .io_a_Z (pippenger_1_pAddPort_1_a_Z[376:0]), //i
    .io_a_T (pippenger_1_pAddPort_1_a_T[376:0]), //i
    .io_b_X (pippenger_1_pAddPort_1_b_X[376:0]), //i
    .io_b_Y (pippenger_1_pAddPort_1_b_Y[376:0]), //i
    .io_b_Z (pippenger_1_pAddPort_1_b_Z[376:0]), //i
    .io_b_T (pippenger_1_pAddPort_1_b_T[376:0]), //i
    .io_s_X (adder_1_io_s_X[376:0]            ), //o
    .io_s_Y (adder_1_io_s_Y[376:0]            ), //o
    .io_s_Z (adder_1_io_s_Z[376:0]            ), //o
    .io_s_T (adder_1_io_s_T[376:0]            ), //o
    .clk    (clk                              ), //i
    .resetn (resetn                           )  //i
  );
  PNeg neg (
    .io_a_X (pippenger_1_pNegPort_a_X[376:0]), //i
    .io_a_Y (pippenger_1_pNegPort_a_Y[376:0]), //i
    .io_a_Z (pippenger_1_pNegPort_a_Z[376:0]), //i
    .io_a_T (pippenger_1_pNegPort_a_T[376:0]), //i
    .io_n_X (neg_io_n_X[376:0]              ), //o
    .io_n_Y (neg_io_n_Y[376:0]              ), //o
    .io_n_Z (neg_io_n_Z[376:0]              ), //o
    .io_n_T (neg_io_n_T[376:0]              ), //o
    .clk    (clk                            ), //i
    .resetn (resetn                         )  //i
  );
  Pippenger pippenger_1 (
    .io_dataIn_valid                (io_dataIn_valid                                                                                     ), //i
    .io_dataIn_ready                (pippenger_1_io_dataIn_ready                                                                         ), //o
    .io_dataIn_payload_last         (io_dataIn_payload_last                                                                              ), //i
    .io_dataIn_payload_fragment_P_X (io_dataIn_payload_fragment_P_X[376:0]                                                               ), //i
    .io_dataIn_payload_fragment_P_Y (io_dataIn_payload_fragment_P_Y[376:0]                                                               ), //i
    .io_dataIn_payload_fragment_P_Z (io_dataIn_payload_fragment_P_Z[376:0]                                                               ), //i
    .io_dataIn_payload_fragment_P_T (io_dataIn_payload_fragment_P_T[376:0]                                                               ), //i
    .io_dataIn_payload_fragment_K   (io_dataIn_payload_fragment_K[252:0]                                                                 ), //i
    .io_dataOut_valid               (pippenger_1_io_dataOut_valid                                                                        ), //o
    .io_dataOut_ready               (io_dataOut_ready                                                                                    ), //i
    .io_dataOut_payload_X           (pippenger_1_io_dataOut_payload_X[376:0]                                                             ), //o
    .io_dataOut_payload_Y           (pippenger_1_io_dataOut_payload_Y[376:0]                                                             ), //o
    .io_dataOut_payload_Z           (pippenger_1_io_dataOut_payload_Z[376:0]                                                             ), //o
    .io_dataOut_payload_T           (pippenger_1_io_dataOut_payload_T[376:0]                                                             ), //o
    .io_pInit_X                     (377'h0                                                                                              ), //i
    .io_pInit_Y                     (377'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001), //i
    .io_pInit_Z                     (377'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001), //i
    .io_pInit_T                     (377'h0                                                                                              ), //i
    .pAddPort_0_a_X                 (pippenger_1_pAddPort_0_a_X[376:0]                                                                   ), //o
    .pAddPort_0_a_Y                 (pippenger_1_pAddPort_0_a_Y[376:0]                                                                   ), //o
    .pAddPort_0_a_Z                 (pippenger_1_pAddPort_0_a_Z[376:0]                                                                   ), //o
    .pAddPort_0_a_T                 (pippenger_1_pAddPort_0_a_T[376:0]                                                                   ), //o
    .pAddPort_0_b_X                 (pippenger_1_pAddPort_0_b_X[376:0]                                                                   ), //o
    .pAddPort_0_b_Y                 (pippenger_1_pAddPort_0_b_Y[376:0]                                                                   ), //o
    .pAddPort_0_b_Z                 (pippenger_1_pAddPort_0_b_Z[376:0]                                                                   ), //o
    .pAddPort_0_b_T                 (pippenger_1_pAddPort_0_b_T[376:0]                                                                   ), //o
    .pAddPort_0_s_X                 (adder_0_io_s_X[376:0]                                                                               ), //i
    .pAddPort_0_s_Y                 (adder_0_io_s_Y[376:0]                                                                               ), //i
    .pAddPort_0_s_Z                 (adder_0_io_s_Z[376:0]                                                                               ), //i
    .pAddPort_0_s_T                 (adder_0_io_s_T[376:0]                                                                               ), //i
    .pAddPort_1_a_X                 (pippenger_1_pAddPort_1_a_X[376:0]                                                                   ), //o
    .pAddPort_1_a_Y                 (pippenger_1_pAddPort_1_a_Y[376:0]                                                                   ), //o
    .pAddPort_1_a_Z                 (pippenger_1_pAddPort_1_a_Z[376:0]                                                                   ), //o
    .pAddPort_1_a_T                 (pippenger_1_pAddPort_1_a_T[376:0]                                                                   ), //o
    .pAddPort_1_b_X                 (pippenger_1_pAddPort_1_b_X[376:0]                                                                   ), //o
    .pAddPort_1_b_Y                 (pippenger_1_pAddPort_1_b_Y[376:0]                                                                   ), //o
    .pAddPort_1_b_Z                 (pippenger_1_pAddPort_1_b_Z[376:0]                                                                   ), //o
    .pAddPort_1_b_T                 (pippenger_1_pAddPort_1_b_T[376:0]                                                                   ), //o
    .pAddPort_1_s_X                 (adder_1_io_s_X[376:0]                                                                               ), //i
    .pAddPort_1_s_Y                 (adder_1_io_s_Y[376:0]                                                                               ), //i
    .pAddPort_1_s_Z                 (adder_1_io_s_Z[376:0]                                                                               ), //i
    .pAddPort_1_s_T                 (adder_1_io_s_T[376:0]                                                                               ), //i
    .pNegPort_a_X                   (pippenger_1_pNegPort_a_X[376:0]                                                                     ), //o
    .pNegPort_a_Y                   (pippenger_1_pNegPort_a_Y[376:0]                                                                     ), //o
    .pNegPort_a_Z                   (pippenger_1_pNegPort_a_Z[376:0]                                                                     ), //o
    .pNegPort_a_T                   (pippenger_1_pNegPort_a_T[376:0]                                                                     ), //o
    .pNegPort_n_X                   (neg_io_n_X[376:0]                                                                                   ), //i
    .pNegPort_n_Y                   (neg_io_n_Y[376:0]                                                                                   ), //i
    .pNegPort_n_Z                   (neg_io_n_Z[376:0]                                                                                   ), //i
    .pNegPort_n_T                   (neg_io_n_T[376:0]                                                                                   ), //i
    .clk                            (clk                                                                                                 ), //i
    .resetn                         (resetn                                                                                              )  //i
  );
  assign io_dataIn_ready = pippenger_1_io_dataIn_ready;
  assign io_dataOut_valid = pippenger_1_io_dataOut_valid;
  assign io_dataOut_payload_X = pippenger_1_io_dataOut_payload_X;
  assign io_dataOut_payload_Y = pippenger_1_io_dataOut_payload_Y;
  assign io_dataOut_payload_Z = pippenger_1_io_dataOut_payload_Z;
  assign io_dataOut_payload_T = pippenger_1_io_dataOut_payload_T;

endmodule

module FIFO (
  input               io_push_valid,
  output              io_push_ready,
  input      [511:0]  io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [511:0]  io_pop_payload,
  output     [7:0]    io_pushPtr,
  output     [7:0]    io_popPtr,
  input               clk,
  input               resetn
);

  reg        [511:0]  _zz_useRam_ram_port1;
  wire       [7:0]    _zz_useRam_pushPtr_valueNext;
  wire       [0:0]    _zz_useRam_pushPtr_valueNext_1;
  wire       [7:0]    _zz_useRam_popPtr_valueNext;
  wire       [0:0]    _zz_useRam_popPtr_valueNext_1;
  wire       [6:0]    _zz_useRam_ram_port;
  wire       [6:0]    _zz_useRam_ram_port_1;
  wire                _zz_useRam_ram_port_2;
  wire       [6:0]    _zz_io_pop_payload_1;
  wire                _zz_io_pop_payload_2;
  reg                 _zz_1;
  reg                 useRam_pushPtr_willIncrement;
  wire                useRam_pushPtr_willClear;
  reg        [7:0]    useRam_pushPtr_valueNext;
  reg        [7:0]    useRam_pushPtr_value;
  reg                 useRam_pushPtr_willOverflowIfInc;
  wire                useRam_pushPtr_willOverflow;
  reg                 useRam_popPtr_willIncrement;
  wire                useRam_popPtr_willClear;
  reg        [7:0]    useRam_popPtr_valueNext;
  reg        [7:0]    useRam_popPtr_value;
  reg                 useRam_popPtr_willOverflowIfInc;
  wire                useRam_popPtr_willOverflow;
  reg                 _zz_io_push_ready;
  wire                io_push_fire;
  reg                 _zz_io_pop_valid;
  wire       [7:0]    _zz_io_pop_payload;
  wire                io_pop_fire;
  reg [511:0] useRam_ram [0:127];

  assign _zz_useRam_pushPtr_valueNext_1 = useRam_pushPtr_willIncrement;
  assign _zz_useRam_pushPtr_valueNext = {7'd0, _zz_useRam_pushPtr_valueNext_1};
  assign _zz_useRam_popPtr_valueNext_1 = useRam_popPtr_willIncrement;
  assign _zz_useRam_popPtr_valueNext = {7'd0, _zz_useRam_popPtr_valueNext_1};
  assign _zz_useRam_ram_port = useRam_pushPtr_value[6:0];
  assign _zz_io_pop_payload_1 = _zz_io_pop_payload[6:0];
  assign _zz_io_pop_payload_2 = 1'b1;
  always @(posedge clk) begin
    if(_zz_1) begin
      useRam_ram[_zz_useRam_ram_port] <= io_push_payload;
    end
  end

  always @(posedge clk) begin
    if(_zz_io_pop_payload_2) begin
      _zz_useRam_ram_port1 <= useRam_ram[_zz_io_pop_payload_1];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    useRam_pushPtr_willIncrement = 1'b0;
    if(io_push_fire) begin
      useRam_pushPtr_willIncrement = 1'b1;
    end
  end

  assign useRam_pushPtr_willClear = 1'b0;
  assign useRam_pushPtr_willOverflow = (useRam_pushPtr_willOverflowIfInc && useRam_pushPtr_willIncrement);
  always @(*) begin
    useRam_pushPtr_valueNext = (useRam_pushPtr_value + _zz_useRam_pushPtr_valueNext);
    if(useRam_pushPtr_willClear) begin
      useRam_pushPtr_valueNext = 8'h0;
    end
  end

  always @(*) begin
    useRam_popPtr_willIncrement = 1'b0;
    if(io_pop_fire) begin
      useRam_popPtr_willIncrement = 1'b1;
    end
  end

  assign useRam_popPtr_willClear = 1'b0;
  assign useRam_popPtr_willOverflow = (useRam_popPtr_willOverflowIfInc && useRam_popPtr_willIncrement);
  always @(*) begin
    useRam_popPtr_valueNext = (useRam_popPtr_value + _zz_useRam_popPtr_valueNext);
    if(useRam_popPtr_willClear) begin
      useRam_popPtr_valueNext = 8'h0;
    end
  end

  assign io_pushPtr = useRam_pushPtr_value;
  assign io_popPtr = useRam_popPtr_value;
  assign io_push_ready = _zz_io_push_ready;
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign io_pop_valid = _zz_io_pop_valid;
  assign _zz_io_pop_payload = useRam_popPtr_valueNext;
  assign io_pop_payload = _zz_useRam_ram_port1;
  assign io_pop_fire = (io_pop_valid && io_pop_ready);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      useRam_pushPtr_value <= 8'h0;
      useRam_pushPtr_willOverflowIfInc <= 1'b0;
      useRam_popPtr_value <= 8'h0;
      useRam_popPtr_willOverflowIfInc <= 1'b0;
      _zz_io_push_ready <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      useRam_pushPtr_value <= useRam_pushPtr_valueNext;
      useRam_pushPtr_willOverflowIfInc <= (useRam_pushPtr_valueNext == 8'hff);
      useRam_popPtr_value <= useRam_popPtr_valueNext;
      useRam_popPtr_willOverflowIfInc <= (useRam_popPtr_valueNext == 8'hff);
      _zz_io_push_ready <= (! ((useRam_pushPtr_valueNext[7] != useRam_popPtr_value[7]) && (useRam_pushPtr_valueNext[6 : 0] == useRam_popPtr_value[6 : 0])));
      _zz_io_pop_valid <= (! (useRam_pushPtr_value == useRam_popPtr_valueNext));
    end
  end


endmodule

module Pippenger (
  input               io_dataIn_valid,
  output              io_dataIn_ready,
  input               io_dataIn_payload_last,
  input      [376:0]  io_dataIn_payload_fragment_P_X,
  input      [376:0]  io_dataIn_payload_fragment_P_Y,
  input      [376:0]  io_dataIn_payload_fragment_P_Z,
  input      [376:0]  io_dataIn_payload_fragment_P_T,
  input      [252:0]  io_dataIn_payload_fragment_K,
  output              io_dataOut_valid,
  input               io_dataOut_ready,
  output     [376:0]  io_dataOut_payload_X,
  output     [376:0]  io_dataOut_payload_Y,
  output     [376:0]  io_dataOut_payload_Z,
  output     [376:0]  io_dataOut_payload_T,
  input      [376:0]  io_pInit_X,
  input      [376:0]  io_pInit_Y,
  input      [376:0]  io_pInit_Z,
  input      [376:0]  io_pInit_T,
  output     [376:0]  pAddPort_0_a_X,
  output     [376:0]  pAddPort_0_a_Y,
  output     [376:0]  pAddPort_0_a_Z,
  output     [376:0]  pAddPort_0_a_T,
  output     [376:0]  pAddPort_0_b_X,
  output     [376:0]  pAddPort_0_b_Y,
  output     [376:0]  pAddPort_0_b_Z,
  output     [376:0]  pAddPort_0_b_T,
  input      [376:0]  pAddPort_0_s_X,
  input      [376:0]  pAddPort_0_s_Y,
  input      [376:0]  pAddPort_0_s_Z,
  input      [376:0]  pAddPort_0_s_T,
  output     [376:0]  pAddPort_1_a_X,
  output     [376:0]  pAddPort_1_a_Y,
  output     [376:0]  pAddPort_1_a_Z,
  output     [376:0]  pAddPort_1_a_T,
  output     [376:0]  pAddPort_1_b_X,
  output     [376:0]  pAddPort_1_b_Y,
  output     [376:0]  pAddPort_1_b_Z,
  output     [376:0]  pAddPort_1_b_T,
  input      [376:0]  pAddPort_1_s_X,
  input      [376:0]  pAddPort_1_s_Y,
  input      [376:0]  pAddPort_1_s_Z,
  input      [376:0]  pAddPort_1_s_T,
  output     [376:0]  pNegPort_a_X,
  output     [376:0]  pNegPort_a_Y,
  output     [376:0]  pNegPort_a_Z,
  output     [376:0]  pNegPort_a_T,
  input      [376:0]  pNegPort_n_X,
  input      [376:0]  pNegPort_n_Y,
  input      [376:0]  pNegPort_n_Z,
  input      [376:0]  pNegPort_n_T,
  input               clk,
  input               resetn
);
  localparam fsm_enumDef_flushing = 5'd1;
  localparam fsm_enumDef_stage1 = 5'd2;
  localparam fsm_enumDef_stage2 = 5'd4;
  localparam fsm_enumDef_stage3 = 5'd8;
  localparam fsm_enumDef_stage3Final = 5'd16;

  reg                 stateRam_0_io_we_0;
  reg                 stateRam_0_io_we_1;
  reg        [15:0]   stateRam_0_io_address_0;
  reg        [15:0]   stateRam_0_io_address_1;
  reg                 stateRam_0_io_flush;
  reg        [15:0]   stateRam_0_io_flushCnt;
  reg                 stateRam_1_1_io_we_0;
  reg                 stateRam_1_1_io_we_1;
  reg        [15:0]   stateRam_1_1_io_address_0;
  reg        [15:0]   stateRam_1_1_io_address_1;
  reg                 stateRam_1_1_io_flush;
  reg        [15:0]   stateRam_1_1_io_flushCnt;
  reg                 dataRam_0_io_we_0;
  reg                 dataRam_0_io_we_1;
  reg        [15:0]   dataRam_0_io_address_0;
  reg        [15:0]   dataRam_0_io_address_1;
  reg        [376:0]  dataRam_0_io_wData_0_X;
  reg        [376:0]  dataRam_0_io_wData_0_Y;
  reg        [376:0]  dataRam_0_io_wData_0_Z;
  reg        [376:0]  dataRam_0_io_wData_0_T;
  reg        [376:0]  dataRam_0_io_wData_1_X;
  reg        [376:0]  dataRam_0_io_wData_1_Y;
  reg        [376:0]  dataRam_0_io_wData_1_Z;
  reg        [376:0]  dataRam_0_io_wData_1_T;
  reg                 dataRam_0_io_state_1;
  reg                 dataRam_1_1_io_we_0;
  reg                 dataRam_1_1_io_we_1;
  reg        [15:0]   dataRam_1_1_io_address_0;
  reg        [15:0]   dataRam_1_1_io_address_1;
  reg        [376:0]  dataRam_1_1_io_wData_0_X;
  reg        [376:0]  dataRam_1_1_io_wData_0_Y;
  reg        [376:0]  dataRam_1_1_io_wData_0_Z;
  reg        [376:0]  dataRam_1_1_io_wData_0_T;
  reg        [376:0]  dataRam_1_1_io_wData_1_X;
  reg        [376:0]  dataRam_1_1_io_wData_1_Y;
  reg        [376:0]  dataRam_1_1_io_wData_1_Z;
  reg        [376:0]  dataRam_1_1_io_wData_1_T;
  reg                 dataRam_1_1_io_state_1;
  reg                 fifo_0_io_dataIn_0_valid;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_a_X;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_a_Y;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_a_Z;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_a_T;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_b_X;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_b_Y;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_b_Z;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_b_T;
  reg        [15:0]   fifo_0_io_dataIn_0_payload_address;
  reg                 fifo_0_io_dataIn_1_valid;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_a_X;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_a_Y;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_a_Z;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_a_T;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_b_X;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_b_Y;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_b_Z;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_b_T;
  reg        [15:0]   fifo_0_io_dataIn_1_payload_address;
  reg                 fifo_1_io_dataIn_0_valid;
  reg        [376:0]  fifo_1_io_dataIn_0_payload_a_X;
  reg        [376:0]  fifo_1_io_dataIn_0_payload_a_Y;
  reg        [376:0]  fifo_1_io_dataIn_0_payload_a_Z;
  reg        [376:0]  fifo_1_io_dataIn_0_payload_a_T;
  reg        [376:0]  fifo_1_io_dataIn_0_payload_b_X;
  reg        [376:0]  fifo_1_io_dataIn_0_payload_b_Y;
  reg        [376:0]  fifo_1_io_dataIn_0_payload_b_Z;
  reg        [376:0]  fifo_1_io_dataIn_0_payload_b_T;
  reg        [15:0]   fifo_1_io_dataIn_0_payload_address;
  reg                 fifo_1_io_dataIn_1_valid;
  reg        [376:0]  fifo_1_io_dataIn_1_payload_a_X;
  reg        [376:0]  fifo_1_io_dataIn_1_payload_a_Y;
  reg        [376:0]  fifo_1_io_dataIn_1_payload_a_Z;
  reg        [376:0]  fifo_1_io_dataIn_1_payload_a_T;
  reg        [376:0]  fifo_1_io_dataIn_1_payload_b_X;
  reg        [376:0]  fifo_1_io_dataIn_1_payload_b_Y;
  reg        [376:0]  fifo_1_io_dataIn_1_payload_b_Z;
  reg        [376:0]  fifo_1_io_dataIn_1_payload_b_T;
  reg        [15:0]   fifo_1_io_dataIn_1_payload_address;
  wire                stateRam_0_io_state_0;
  wire                stateRam_0_io_state_1;
  wire                stateRam_1_1_io_state_0;
  wire                stateRam_1_1_io_state_1;
  wire       [376:0]  dataRam_0_io_rData_0_X;
  wire       [376:0]  dataRam_0_io_rData_0_Y;
  wire       [376:0]  dataRam_0_io_rData_0_Z;
  wire       [376:0]  dataRam_0_io_rData_0_T;
  wire       [376:0]  dataRam_0_io_rData_1_X;
  wire       [376:0]  dataRam_0_io_rData_1_Y;
  wire       [376:0]  dataRam_0_io_rData_1_Z;
  wire       [376:0]  dataRam_0_io_rData_1_T;
  wire       [376:0]  dataRam_1_1_io_rData_0_X;
  wire       [376:0]  dataRam_1_1_io_rData_0_Y;
  wire       [376:0]  dataRam_1_1_io_rData_0_Z;
  wire       [376:0]  dataRam_1_1_io_rData_0_T;
  wire       [376:0]  dataRam_1_1_io_rData_1_X;
  wire       [376:0]  dataRam_1_1_io_rData_1_Y;
  wire       [376:0]  dataRam_1_1_io_rData_1_Z;
  wire       [376:0]  dataRam_1_1_io_rData_1_T;
  wire                fifo_0_io_dataOut_valid;
  wire       [376:0]  fifo_0_io_dataOut_payload_a_X;
  wire       [376:0]  fifo_0_io_dataOut_payload_a_Y;
  wire       [376:0]  fifo_0_io_dataOut_payload_a_Z;
  wire       [376:0]  fifo_0_io_dataOut_payload_a_T;
  wire       [376:0]  fifo_0_io_dataOut_payload_b_X;
  wire       [376:0]  fifo_0_io_dataOut_payload_b_Y;
  wire       [376:0]  fifo_0_io_dataOut_payload_b_Z;
  wire       [376:0]  fifo_0_io_dataOut_payload_b_T;
  wire       [15:0]   fifo_0_io_dataOut_payload_address;
  wire                fifo_1_io_dataOut_valid;
  wire       [376:0]  fifo_1_io_dataOut_payload_a_X;
  wire       [376:0]  fifo_1_io_dataOut_payload_a_Y;
  wire       [376:0]  fifo_1_io_dataOut_payload_a_Z;
  wire       [376:0]  fifo_1_io_dataOut_payload_a_T;
  wire       [376:0]  fifo_1_io_dataOut_payload_b_X;
  wire       [376:0]  fifo_1_io_dataOut_payload_b_Y;
  wire       [376:0]  fifo_1_io_dataOut_payload_b_Z;
  wire       [376:0]  fifo_1_io_dataOut_payload_b_T;
  wire       [15:0]   fifo_1_io_dataOut_payload_address;
  wire       [226:0]  _zz_dataInBuffer_dataReg_fragment_K;
  wire       [15:0]   _zz_flushing_flushCnt_valueNext;
  wire       [0:0]    _zz_flushing_flushCnt_valueNext_1;
  wire       [31:0]   _zz_stage1_NCnt_valueNext;
  wire       [0:0]    _zz_stage1_NCnt_valueNext_1;
  wire       [3:0]    _zz_stage1_GCnt_valueNext;
  wire       [0:0]    _zz_stage1_GCnt_valueNext_1;
  wire       [8:0]    _zz_stage1_emptyCnt_valueNext;
  wire       [0:0]    _zz_stage1_emptyCnt_valueNext_1;
  wire       [13:0]   _zz_stage1_inputBarrelID_0_1;
  wire       [1:0]    _zz_stage1_inputBarrelID_0_2;
  wire       [13:0]   _zz_stage1_inputBarrelID_1;
  wire       [1:0]    _zz_stage1_inputBarrelID_1_1;
  wire       [12:0]   _zz__zz_stage1_inputBarrelIDAbs_0;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0_1;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0_2;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0_3;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0_4;
  wire       [0:0]    _zz_stage1_inputBarrelIDAbs_0_5;
  wire       [12:0]   _zz__zz_stage1_inputBarrelIDAbs_1;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_1_1;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_1_2;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_1_3;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_1_4;
  wire       [0:0]    _zz_stage1_inputBarrelIDAbs_1_5;
  wire       [12:0]   _zz__zz_stage1_inputValid_0;
  wire       [12:0]   _zz__zz_stage1_inputValid_1;
  wire       [11:0]   _zz_stage2_wCnt_valueNext;
  wire       [0:0]    _zz_stage2_wCnt_valueNext_1;
  wire       [3:0]    _zz_stage2_GCnt_valueNext;
  wire       [0:0]    _zz_stage2_GCnt_valueNext_1;
  wire       [1:0]    _zz_stage2_calCnt_valueNext;
  wire       [0:0]    _zz_stage2_calCnt_valueNext_1;
  wire       [8:0]    _zz_stage2_waitCnt_valueNext;
  wire       [0:0]    _zz_stage2_waitCnt_valueNext_1;
  wire       [3:0]    _zz_stage3_GCnt_valueNext;
  wire       [0:0]    _zz_stage3_GCnt_valueNext_1;
  wire       [4:0]    _zz_stage3_doubleCnt_valueNext;
  wire       [0:0]    _zz_stage3_doubleCnt_valueNext_1;
  wire       [8:0]    _zz_stage3_doubleWaitCnt_valueNext;
  wire       [0:0]    _zz_stage3_doubleWaitCnt_valueNext_1;
  wire       [8:0]    _zz_stage3_addWaitCnt_valueNext;
  wire       [0:0]    _zz_stage3_addWaitCnt_valueNext_1;
  wire       [3:0]    _zz_stage3Final_doubleCnt_valueNext;
  wire       [0:0]    _zz_stage3Final_doubleCnt_valueNext_1;
  wire       [8:0]    _zz_stage3Final_doubleWaitCnt_valueNext;
  wire       [0:0]    _zz_stage3Final_doubleWaitCnt_valueNext_1;
  wire       [8:0]    _zz_stage3Final_addWaitCnt_valueNext;
  wire       [0:0]    _zz_stage3Final_addWaitCnt_valueNext_1;
  wire       [11:0]   _zz_io_address_0;
  wire       [11:0]   _zz_io_address_0_1;
  wire       [11:0]   _zz_io_address_0_2;
  wire       [11:0]   _zz_io_address_1;
  wire       [11:0]   _zz_io_address_1_1;
  wire       [11:0]   _zz_io_address_1_2;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address_1;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address_2;
  wire       [11:0]   _zz_io_address_0_3;
  wire       [11:0]   _zz_io_address_0_4;
  wire       [11:0]   _zz_io_address_0_5;
  wire       [11:0]   _zz_io_address_1_3;
  wire       [11:0]   _zz_io_address_1_4;
  wire       [11:0]   _zz_io_address_1_5;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address_30;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address_30_1;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address_30_2;
  wire       [3:0]    _zz_io_address_1_6;
  wire       [3:0]    _zz_io_address_1_7;
  wire       [0:0]    _zz_io_address_1_8;
  wire       [3:0]    _zz__zz_io_dataIn_1_payload_address_60;
  wire       [0:0]    _zz__zz_io_dataIn_1_payload_address_60_1;
  wire       [3:0]    _zz_io_address_1_9;
  wire       [3:0]    _zz_io_address_1_10;
  wire       [0:0]    _zz_io_address_1_11;
  wire       [3:0]    _zz__zz_io_dataIn_1_payload_address_90;
  wire       [0:0]    _zz__zz_io_dataIn_1_payload_address_90_1;
  wire                dataInBuffer_bufferOut_valid;
  reg                 dataInBuffer_bufferOut_ready;
  wire                dataInBuffer_bufferOut_payload_last;
  wire       [376:0]  dataInBuffer_bufferOut_payload_fragment_P_X;
  wire       [376:0]  dataInBuffer_bufferOut_payload_fragment_P_Y;
  wire       [376:0]  dataInBuffer_bufferOut_payload_fragment_P_Z;
  wire       [376:0]  dataInBuffer_bufferOut_payload_fragment_P_T;
  wire       [252:0]  dataInBuffer_bufferOut_payload_fragment_K;
  reg                 dataInBuffer_shift;
  reg                 dataInBuffer_validReg;
  reg                 dataInBuffer_dataReg_last;
  reg        [376:0]  dataInBuffer_dataReg_fragment_P_X;
  reg        [376:0]  dataInBuffer_dataReg_fragment_P_Y;
  reg        [376:0]  dataInBuffer_dataReg_fragment_P_Z;
  reg        [376:0]  dataInBuffer_dataReg_fragment_P_T;
  reg        [252:0]  dataInBuffer_dataReg_fragment_K;
  wire                shiftRegs_validIn_0;
  wire                shiftRegs_validIn_1;
  wire       [15:0]   shiftRegs_addressIn_0;
  wire       [15:0]   shiftRegs_addressIn_1;
  reg                 shiftRegs_validIn_delay_1_0;
  reg                 shiftRegs_validIn_delay_1_1;
  reg                 shiftRegs_validIn_delay_2_0;
  reg                 shiftRegs_validIn_delay_2_1;
  reg                 shiftRegs_validIn_delay_3_0;
  reg                 shiftRegs_validIn_delay_3_1;
  reg                 shiftRegs_validIn_delay_4_0;
  reg                 shiftRegs_validIn_delay_4_1;
  reg                 shiftRegs_validIn_delay_5_0;
  reg                 shiftRegs_validIn_delay_5_1;
  reg                 shiftRegs_validIn_delay_6_0;
  reg                 shiftRegs_validIn_delay_6_1;
  reg                 shiftRegs_validIn_delay_7_0;
  reg                 shiftRegs_validIn_delay_7_1;
  reg                 shiftRegs_validIn_delay_8_0;
  reg                 shiftRegs_validIn_delay_8_1;
  reg                 shiftRegs_validIn_delay_9_0;
  reg                 shiftRegs_validIn_delay_9_1;
  reg                 shiftRegs_validIn_delay_10_0;
  reg                 shiftRegs_validIn_delay_10_1;
  reg                 shiftRegs_validIn_delay_11_0;
  reg                 shiftRegs_validIn_delay_11_1;
  reg                 shiftRegs_validIn_delay_12_0;
  reg                 shiftRegs_validIn_delay_12_1;
  reg                 shiftRegs_validIn_delay_13_0;
  reg                 shiftRegs_validIn_delay_13_1;
  reg                 shiftRegs_validIn_delay_14_0;
  reg                 shiftRegs_validIn_delay_14_1;
  reg                 shiftRegs_validIn_delay_15_0;
  reg                 shiftRegs_validIn_delay_15_1;
  reg                 shiftRegs_validIn_delay_16_0;
  reg                 shiftRegs_validIn_delay_16_1;
  reg                 shiftRegs_validIn_delay_17_0;
  reg                 shiftRegs_validIn_delay_17_1;
  reg                 shiftRegs_validIn_delay_18_0;
  reg                 shiftRegs_validIn_delay_18_1;
  reg                 shiftRegs_validIn_delay_19_0;
  reg                 shiftRegs_validIn_delay_19_1;
  reg                 shiftRegs_validIn_delay_20_0;
  reg                 shiftRegs_validIn_delay_20_1;
  reg                 shiftRegs_validIn_delay_21_0;
  reg                 shiftRegs_validIn_delay_21_1;
  reg                 shiftRegs_validIn_delay_22_0;
  reg                 shiftRegs_validIn_delay_22_1;
  reg                 shiftRegs_validIn_delay_23_0;
  reg                 shiftRegs_validIn_delay_23_1;
  reg                 shiftRegs_validIn_delay_24_0;
  reg                 shiftRegs_validIn_delay_24_1;
  reg                 shiftRegs_validIn_delay_25_0;
  reg                 shiftRegs_validIn_delay_25_1;
  reg                 shiftRegs_validIn_delay_26_0;
  reg                 shiftRegs_validIn_delay_26_1;
  reg                 shiftRegs_validIn_delay_27_0;
  reg                 shiftRegs_validIn_delay_27_1;
  reg                 shiftRegs_validIn_delay_28_0;
  reg                 shiftRegs_validIn_delay_28_1;
  reg                 shiftRegs_validIn_delay_29_0;
  reg                 shiftRegs_validIn_delay_29_1;
  reg                 shiftRegs_validIn_delay_30_0;
  reg                 shiftRegs_validIn_delay_30_1;
  reg                 shiftRegs_validIn_delay_31_0;
  reg                 shiftRegs_validIn_delay_31_1;
  reg                 shiftRegs_validIn_delay_32_0;
  reg                 shiftRegs_validIn_delay_32_1;
  reg                 shiftRegs_validIn_delay_33_0;
  reg                 shiftRegs_validIn_delay_33_1;
  reg                 shiftRegs_validIn_delay_34_0;
  reg                 shiftRegs_validIn_delay_34_1;
  reg                 shiftRegs_validIn_delay_35_0;
  reg                 shiftRegs_validIn_delay_35_1;
  reg                 shiftRegs_validIn_delay_36_0;
  reg                 shiftRegs_validIn_delay_36_1;
  reg                 shiftRegs_validIn_delay_37_0;
  reg                 shiftRegs_validIn_delay_37_1;
  reg                 shiftRegs_validIn_delay_38_0;
  reg                 shiftRegs_validIn_delay_38_1;
  reg                 shiftRegs_validIn_delay_39_0;
  reg                 shiftRegs_validIn_delay_39_1;
  reg                 shiftRegs_validIn_delay_40_0;
  reg                 shiftRegs_validIn_delay_40_1;
  reg                 shiftRegs_validIn_delay_41_0;
  reg                 shiftRegs_validIn_delay_41_1;
  reg                 shiftRegs_validIn_delay_42_0;
  reg                 shiftRegs_validIn_delay_42_1;
  reg                 shiftRegs_validIn_delay_43_0;
  reg                 shiftRegs_validIn_delay_43_1;
  reg                 shiftRegs_validIn_delay_44_0;
  reg                 shiftRegs_validIn_delay_44_1;
  reg                 shiftRegs_validIn_delay_45_0;
  reg                 shiftRegs_validIn_delay_45_1;
  reg                 shiftRegs_validIn_delay_46_0;
  reg                 shiftRegs_validIn_delay_46_1;
  reg                 shiftRegs_validIn_delay_47_0;
  reg                 shiftRegs_validIn_delay_47_1;
  reg                 shiftRegs_validIn_delay_48_0;
  reg                 shiftRegs_validIn_delay_48_1;
  reg                 shiftRegs_validIn_delay_49_0;
  reg                 shiftRegs_validIn_delay_49_1;
  reg                 shiftRegs_validIn_delay_50_0;
  reg                 shiftRegs_validIn_delay_50_1;
  reg                 shiftRegs_validIn_delay_51_0;
  reg                 shiftRegs_validIn_delay_51_1;
  reg                 shiftRegs_validIn_delay_52_0;
  reg                 shiftRegs_validIn_delay_52_1;
  reg                 shiftRegs_validIn_delay_53_0;
  reg                 shiftRegs_validIn_delay_53_1;
  reg                 shiftRegs_validIn_delay_54_0;
  reg                 shiftRegs_validIn_delay_54_1;
  reg                 shiftRegs_validIn_delay_55_0;
  reg                 shiftRegs_validIn_delay_55_1;
  reg                 shiftRegs_validIn_delay_56_0;
  reg                 shiftRegs_validIn_delay_56_1;
  reg                 shiftRegs_validIn_delay_57_0;
  reg                 shiftRegs_validIn_delay_57_1;
  reg                 shiftRegs_validIn_delay_58_0;
  reg                 shiftRegs_validIn_delay_58_1;
  reg                 shiftRegs_validIn_delay_59_0;
  reg                 shiftRegs_validIn_delay_59_1;
  reg                 shiftRegs_validIn_delay_60_0;
  reg                 shiftRegs_validIn_delay_60_1;
  reg                 shiftRegs_validIn_delay_61_0;
  reg                 shiftRegs_validIn_delay_61_1;
  reg                 shiftRegs_validIn_delay_62_0;
  reg                 shiftRegs_validIn_delay_62_1;
  reg                 shiftRegs_validIn_delay_63_0;
  reg                 shiftRegs_validIn_delay_63_1;
  reg                 shiftRegs_validIn_delay_64_0;
  reg                 shiftRegs_validIn_delay_64_1;
  reg                 shiftRegs_validIn_delay_65_0;
  reg                 shiftRegs_validIn_delay_65_1;
  reg                 shiftRegs_validIn_delay_66_0;
  reg                 shiftRegs_validIn_delay_66_1;
  reg                 shiftRegs_validIn_delay_67_0;
  reg                 shiftRegs_validIn_delay_67_1;
  reg                 shiftRegs_validIn_delay_68_0;
  reg                 shiftRegs_validIn_delay_68_1;
  reg                 shiftRegs_validIn_delay_69_0;
  reg                 shiftRegs_validIn_delay_69_1;
  reg                 shiftRegs_validIn_delay_70_0;
  reg                 shiftRegs_validIn_delay_70_1;
  reg                 shiftRegs_validIn_delay_71_0;
  reg                 shiftRegs_validIn_delay_71_1;
  reg                 shiftRegs_validIn_delay_72_0;
  reg                 shiftRegs_validIn_delay_72_1;
  reg                 shiftRegs_validIn_delay_73_0;
  reg                 shiftRegs_validIn_delay_73_1;
  reg                 shiftRegs_validIn_delay_74_0;
  reg                 shiftRegs_validIn_delay_74_1;
  reg                 shiftRegs_validIn_delay_75_0;
  reg                 shiftRegs_validIn_delay_75_1;
  reg                 shiftRegs_validIn_delay_76_0;
  reg                 shiftRegs_validIn_delay_76_1;
  reg                 shiftRegs_validIn_delay_77_0;
  reg                 shiftRegs_validIn_delay_77_1;
  reg                 shiftRegs_validIn_delay_78_0;
  reg                 shiftRegs_validIn_delay_78_1;
  reg                 shiftRegs_validIn_delay_79_0;
  reg                 shiftRegs_validIn_delay_79_1;
  reg                 shiftRegs_validIn_delay_80_0;
  reg                 shiftRegs_validIn_delay_80_1;
  reg                 shiftRegs_validIn_delay_81_0;
  reg                 shiftRegs_validIn_delay_81_1;
  reg                 shiftRegs_validIn_delay_82_0;
  reg                 shiftRegs_validIn_delay_82_1;
  reg                 shiftRegs_validIn_delay_83_0;
  reg                 shiftRegs_validIn_delay_83_1;
  reg                 shiftRegs_validIn_delay_84_0;
  reg                 shiftRegs_validIn_delay_84_1;
  reg                 shiftRegs_validIn_delay_85_0;
  reg                 shiftRegs_validIn_delay_85_1;
  reg                 shiftRegs_validIn_delay_86_0;
  reg                 shiftRegs_validIn_delay_86_1;
  reg                 shiftRegs_validIn_delay_87_0;
  reg                 shiftRegs_validIn_delay_87_1;
  reg                 shiftRegs_validIn_delay_88_0;
  reg                 shiftRegs_validIn_delay_88_1;
  reg                 shiftRegs_validIn_delay_89_0;
  reg                 shiftRegs_validIn_delay_89_1;
  reg                 shiftRegs_validIn_delay_90_0;
  reg                 shiftRegs_validIn_delay_90_1;
  reg                 shiftRegs_validIn_delay_91_0;
  reg                 shiftRegs_validIn_delay_91_1;
  reg                 shiftRegs_validIn_delay_92_0;
  reg                 shiftRegs_validIn_delay_92_1;
  reg                 shiftRegs_validIn_delay_93_0;
  reg                 shiftRegs_validIn_delay_93_1;
  reg                 shiftRegs_validIn_delay_94_0;
  reg                 shiftRegs_validIn_delay_94_1;
  reg                 shiftRegs_validIn_delay_95_0;
  reg                 shiftRegs_validIn_delay_95_1;
  reg                 shiftRegs_validIn_delay_96_0;
  reg                 shiftRegs_validIn_delay_96_1;
  reg                 shiftRegs_validIn_delay_97_0;
  reg                 shiftRegs_validIn_delay_97_1;
  reg                 shiftRegs_validIn_delay_98_0;
  reg                 shiftRegs_validIn_delay_98_1;
  reg                 shiftRegs_validIn_delay_99_0;
  reg                 shiftRegs_validIn_delay_99_1;
  reg                 shiftRegs_validIn_delay_100_0;
  reg                 shiftRegs_validIn_delay_100_1;
  reg                 shiftRegs_validIn_delay_101_0;
  reg                 shiftRegs_validIn_delay_101_1;
  reg                 shiftRegs_validIn_delay_102_0;
  reg                 shiftRegs_validIn_delay_102_1;
  reg                 shiftRegs_validIn_delay_103_0;
  reg                 shiftRegs_validIn_delay_103_1;
  reg                 shiftRegs_validIn_delay_104_0;
  reg                 shiftRegs_validIn_delay_104_1;
  reg                 shiftRegs_validIn_delay_105_0;
  reg                 shiftRegs_validIn_delay_105_1;
  reg                 shiftRegs_validIn_delay_106_0;
  reg                 shiftRegs_validIn_delay_106_1;
  reg                 shiftRegs_validIn_delay_107_0;
  reg                 shiftRegs_validIn_delay_107_1;
  reg                 shiftRegs_validIn_delay_108_0;
  reg                 shiftRegs_validIn_delay_108_1;
  reg                 shiftRegs_validIn_delay_109_0;
  reg                 shiftRegs_validIn_delay_109_1;
  reg                 shiftRegs_validIn_delay_110_0;
  reg                 shiftRegs_validIn_delay_110_1;
  reg                 shiftRegs_validIn_delay_111_0;
  reg                 shiftRegs_validIn_delay_111_1;
  reg                 shiftRegs_validIn_delay_112_0;
  reg                 shiftRegs_validIn_delay_112_1;
  reg                 shiftRegs_validIn_delay_113_0;
  reg                 shiftRegs_validIn_delay_113_1;
  reg                 shiftRegs_validIn_delay_114_0;
  reg                 shiftRegs_validIn_delay_114_1;
  reg                 shiftRegs_validIn_delay_115_0;
  reg                 shiftRegs_validIn_delay_115_1;
  reg                 shiftRegs_validIn_delay_116_0;
  reg                 shiftRegs_validIn_delay_116_1;
  reg                 shiftRegs_validIn_delay_117_0;
  reg                 shiftRegs_validIn_delay_117_1;
  reg                 shiftRegs_validIn_delay_118_0;
  reg                 shiftRegs_validIn_delay_118_1;
  reg                 shiftRegs_validIn_delay_119_0;
  reg                 shiftRegs_validIn_delay_119_1;
  reg                 shiftRegs_validIn_delay_120_0;
  reg                 shiftRegs_validIn_delay_120_1;
  reg                 shiftRegs_validIn_delay_121_0;
  reg                 shiftRegs_validIn_delay_121_1;
  reg                 shiftRegs_validIn_delay_122_0;
  reg                 shiftRegs_validIn_delay_122_1;
  reg                 shiftRegs_validIn_delay_123_0;
  reg                 shiftRegs_validIn_delay_123_1;
  reg                 shiftRegs_validIn_delay_124_0;
  reg                 shiftRegs_validIn_delay_124_1;
  reg                 shiftRegs_validIn_delay_125_0;
  reg                 shiftRegs_validIn_delay_125_1;
  reg                 shiftRegs_validIn_delay_126_0;
  reg                 shiftRegs_validIn_delay_126_1;
  reg                 shiftRegs_validIn_delay_127_0;
  reg                 shiftRegs_validIn_delay_127_1;
  reg                 shiftRegs_validIn_delay_128_0;
  reg                 shiftRegs_validIn_delay_128_1;
  reg                 shiftRegs_validIn_delay_129_0;
  reg                 shiftRegs_validIn_delay_129_1;
  reg                 shiftRegs_validIn_delay_130_0;
  reg                 shiftRegs_validIn_delay_130_1;
  reg                 shiftRegs_validIn_delay_131_0;
  reg                 shiftRegs_validIn_delay_131_1;
  reg                 shiftRegs_validIn_delay_132_0;
  reg                 shiftRegs_validIn_delay_132_1;
  reg                 shiftRegs_validIn_delay_133_0;
  reg                 shiftRegs_validIn_delay_133_1;
  reg                 shiftRegs_validIn_delay_134_0;
  reg                 shiftRegs_validIn_delay_134_1;
  reg                 shiftRegs_validIn_delay_135_0;
  reg                 shiftRegs_validIn_delay_135_1;
  reg                 shiftRegs_validIn_delay_136_0;
  reg                 shiftRegs_validIn_delay_136_1;
  reg                 shiftRegs_validIn_delay_137_0;
  reg                 shiftRegs_validIn_delay_137_1;
  reg                 shiftRegs_validIn_delay_138_0;
  reg                 shiftRegs_validIn_delay_138_1;
  reg                 shiftRegs_validIn_delay_139_0;
  reg                 shiftRegs_validIn_delay_139_1;
  reg                 shiftRegs_validIn_delay_140_0;
  reg                 shiftRegs_validIn_delay_140_1;
  reg                 shiftRegs_validIn_delay_141_0;
  reg                 shiftRegs_validIn_delay_141_1;
  reg                 shiftRegs_validIn_delay_142_0;
  reg                 shiftRegs_validIn_delay_142_1;
  reg                 shiftRegs_validIn_delay_143_0;
  reg                 shiftRegs_validIn_delay_143_1;
  reg                 shiftRegs_validIn_delay_144_0;
  reg                 shiftRegs_validIn_delay_144_1;
  reg                 shiftRegs_validIn_delay_145_0;
  reg                 shiftRegs_validIn_delay_145_1;
  reg                 shiftRegs_validIn_delay_146_0;
  reg                 shiftRegs_validIn_delay_146_1;
  reg                 shiftRegs_validIn_delay_147_0;
  reg                 shiftRegs_validIn_delay_147_1;
  reg                 shiftRegs_validIn_delay_148_0;
  reg                 shiftRegs_validIn_delay_148_1;
  reg                 shiftRegs_validIn_delay_149_0;
  reg                 shiftRegs_validIn_delay_149_1;
  reg                 shiftRegs_validIn_delay_150_0;
  reg                 shiftRegs_validIn_delay_150_1;
  reg                 shiftRegs_validIn_delay_151_0;
  reg                 shiftRegs_validIn_delay_151_1;
  reg                 shiftRegs_validIn_delay_152_0;
  reg                 shiftRegs_validIn_delay_152_1;
  reg                 shiftRegs_validIn_delay_153_0;
  reg                 shiftRegs_validIn_delay_153_1;
  reg                 shiftRegs_validIn_delay_154_0;
  reg                 shiftRegs_validIn_delay_154_1;
  reg                 shiftRegs_validIn_delay_155_0;
  reg                 shiftRegs_validIn_delay_155_1;
  reg                 shiftRegs_validIn_delay_156_0;
  reg                 shiftRegs_validIn_delay_156_1;
  reg                 shiftRegs_validIn_delay_157_0;
  reg                 shiftRegs_validIn_delay_157_1;
  reg                 shiftRegs_validIn_delay_158_0;
  reg                 shiftRegs_validIn_delay_158_1;
  reg                 shiftRegs_validIn_delay_159_0;
  reg                 shiftRegs_validIn_delay_159_1;
  reg                 shiftRegs_validIn_delay_160_0;
  reg                 shiftRegs_validIn_delay_160_1;
  reg                 shiftRegs_validIn_delay_161_0;
  reg                 shiftRegs_validIn_delay_161_1;
  reg                 shiftRegs_validIn_delay_162_0;
  reg                 shiftRegs_validIn_delay_162_1;
  reg                 shiftRegs_validIn_delay_163_0;
  reg                 shiftRegs_validIn_delay_163_1;
  reg                 shiftRegs_validIn_delay_164_0;
  reg                 shiftRegs_validIn_delay_164_1;
  reg                 shiftRegs_validIn_delay_165_0;
  reg                 shiftRegs_validIn_delay_165_1;
  reg                 shiftRegs_validIn_delay_166_0;
  reg                 shiftRegs_validIn_delay_166_1;
  reg                 shiftRegs_validIn_delay_167_0;
  reg                 shiftRegs_validIn_delay_167_1;
  reg                 shiftRegs_validIn_delay_168_0;
  reg                 shiftRegs_validIn_delay_168_1;
  reg                 shiftRegs_validIn_delay_169_0;
  reg                 shiftRegs_validIn_delay_169_1;
  reg                 shiftRegs_validIn_delay_170_0;
  reg                 shiftRegs_validIn_delay_170_1;
  reg                 shiftRegs_validIn_delay_171_0;
  reg                 shiftRegs_validIn_delay_171_1;
  reg                 shiftRegs_validIn_delay_172_0;
  reg                 shiftRegs_validIn_delay_172_1;
  reg                 shiftRegs_validIn_delay_173_0;
  reg                 shiftRegs_validIn_delay_173_1;
  reg                 shiftRegs_validIn_delay_174_0;
  reg                 shiftRegs_validIn_delay_174_1;
  reg                 shiftRegs_validIn_delay_175_0;
  reg                 shiftRegs_validIn_delay_175_1;
  reg                 shiftRegs_validIn_delay_176_0;
  reg                 shiftRegs_validIn_delay_176_1;
  reg                 shiftRegs_validIn_delay_177_0;
  reg                 shiftRegs_validIn_delay_177_1;
  reg                 shiftRegs_validIn_delay_178_0;
  reg                 shiftRegs_validIn_delay_178_1;
  reg                 shiftRegs_validIn_delay_179_0;
  reg                 shiftRegs_validIn_delay_179_1;
  reg                 shiftRegs_validIn_delay_180_0;
  reg                 shiftRegs_validIn_delay_180_1;
  reg                 shiftRegs_validIn_delay_181_0;
  reg                 shiftRegs_validIn_delay_181_1;
  reg                 shiftRegs_validIn_delay_182_0;
  reg                 shiftRegs_validIn_delay_182_1;
  reg                 shiftRegs_validIn_delay_183_0;
  reg                 shiftRegs_validIn_delay_183_1;
  reg                 shiftRegs_validIn_delay_184_0;
  reg                 shiftRegs_validIn_delay_184_1;
  reg                 shiftRegs_validIn_delay_185_0;
  reg                 shiftRegs_validIn_delay_185_1;
  reg                 shiftRegs_validIn_delay_186_0;
  reg                 shiftRegs_validIn_delay_186_1;
  reg                 shiftRegs_validIn_delay_187_0;
  reg                 shiftRegs_validIn_delay_187_1;
  reg                 shiftRegs_validIn_delay_188_0;
  reg                 shiftRegs_validIn_delay_188_1;
  reg                 shiftRegs_validIn_delay_189_0;
  reg                 shiftRegs_validIn_delay_189_1;
  reg                 shiftRegs_validIn_delay_190_0;
  reg                 shiftRegs_validIn_delay_190_1;
  reg                 shiftRegs_validIn_delay_191_0;
  reg                 shiftRegs_validIn_delay_191_1;
  reg                 shiftRegs_validIn_delay_192_0;
  reg                 shiftRegs_validIn_delay_192_1;
  reg                 shiftRegs_validIn_delay_193_0;
  reg                 shiftRegs_validIn_delay_193_1;
  reg                 shiftRegs_validIn_delay_194_0;
  reg                 shiftRegs_validIn_delay_194_1;
  reg                 shiftRegs_validIn_delay_195_0;
  reg                 shiftRegs_validIn_delay_195_1;
  reg                 shiftRegs_validIn_delay_196_0;
  reg                 shiftRegs_validIn_delay_196_1;
  reg                 shiftRegs_validIn_delay_197_0;
  reg                 shiftRegs_validIn_delay_197_1;
  reg                 shiftRegs_validIn_delay_198_0;
  reg                 shiftRegs_validIn_delay_198_1;
  reg                 shiftRegs_validIn_delay_199_0;
  reg                 shiftRegs_validIn_delay_199_1;
  reg                 shiftRegs_validIn_delay_200_0;
  reg                 shiftRegs_validIn_delay_200_1;
  reg                 shiftRegs_validIn_delay_201_0;
  reg                 shiftRegs_validIn_delay_201_1;
  reg                 shiftRegs_validIn_delay_202_0;
  reg                 shiftRegs_validIn_delay_202_1;
  reg                 shiftRegs_validIn_delay_203_0;
  reg                 shiftRegs_validIn_delay_203_1;
  reg                 shiftRegs_validIn_delay_204_0;
  reg                 shiftRegs_validIn_delay_204_1;
  reg                 shiftRegs_validIn_delay_205_0;
  reg                 shiftRegs_validIn_delay_205_1;
  reg                 shiftRegs_validIn_delay_206_0;
  reg                 shiftRegs_validIn_delay_206_1;
  reg                 shiftRegs_validIn_delay_207_0;
  reg                 shiftRegs_validIn_delay_207_1;
  reg                 shiftRegs_validIn_delay_208_0;
  reg                 shiftRegs_validIn_delay_208_1;
  reg                 shiftRegs_validIn_delay_209_0;
  reg                 shiftRegs_validIn_delay_209_1;
  reg                 shiftRegs_validIn_delay_210_0;
  reg                 shiftRegs_validIn_delay_210_1;
  reg                 shiftRegs_validIn_delay_211_0;
  reg                 shiftRegs_validIn_delay_211_1;
  reg                 shiftRegs_validIn_delay_212_0;
  reg                 shiftRegs_validIn_delay_212_1;
  reg                 shiftRegs_validIn_delay_213_0;
  reg                 shiftRegs_validIn_delay_213_1;
  reg                 shiftRegs_validIn_delay_214_0;
  reg                 shiftRegs_validIn_delay_214_1;
  reg                 shiftRegs_validIn_delay_215_0;
  reg                 shiftRegs_validIn_delay_215_1;
  reg                 shiftRegs_validIn_delay_216_0;
  reg                 shiftRegs_validIn_delay_216_1;
  reg                 shiftRegs_validIn_delay_217_0;
  reg                 shiftRegs_validIn_delay_217_1;
  reg                 shiftRegs_validIn_delay_218_0;
  reg                 shiftRegs_validIn_delay_218_1;
  reg                 shiftRegs_validIn_delay_219_0;
  reg                 shiftRegs_validIn_delay_219_1;
  reg                 shiftRegs_validIn_delay_220_0;
  reg                 shiftRegs_validIn_delay_220_1;
  reg                 shiftRegs_validIn_delay_221_0;
  reg                 shiftRegs_validIn_delay_221_1;
  reg                 shiftRegs_validIn_delay_222_0;
  reg                 shiftRegs_validIn_delay_222_1;
  reg                 shiftRegs_validIn_delay_223_0;
  reg                 shiftRegs_validIn_delay_223_1;
  reg                 shiftRegs_validIn_delay_224_0;
  reg                 shiftRegs_validIn_delay_224_1;
  reg                 shiftRegs_validIn_delay_225_0;
  reg                 shiftRegs_validIn_delay_225_1;
  reg                 shiftRegs_validIn_delay_226_0;
  reg                 shiftRegs_validIn_delay_226_1;
  reg                 shiftRegs_validIn_delay_227_0;
  reg                 shiftRegs_validIn_delay_227_1;
  reg                 shiftRegs_validIn_delay_228_0;
  reg                 shiftRegs_validIn_delay_228_1;
  reg                 shiftRegs_validIn_delay_229_0;
  reg                 shiftRegs_validIn_delay_229_1;
  reg                 shiftRegs_validIn_delay_230_0;
  reg                 shiftRegs_validIn_delay_230_1;
  reg                 shiftRegs_validIn_delay_231_0;
  reg                 shiftRegs_validIn_delay_231_1;
  reg                 shiftRegs_validIn_delay_232_0;
  reg                 shiftRegs_validIn_delay_232_1;
  reg                 shiftRegs_validIn_delay_233_0;
  reg                 shiftRegs_validIn_delay_233_1;
  reg                 shiftRegs_validIn_delay_234_0;
  reg                 shiftRegs_validIn_delay_234_1;
  reg                 shiftRegs_validIn_delay_235_0;
  reg                 shiftRegs_validIn_delay_235_1;
  reg                 shiftRegs_validIn_delay_236_0;
  reg                 shiftRegs_validIn_delay_236_1;
  reg                 shiftRegs_validIn_delay_237_0;
  reg                 shiftRegs_validIn_delay_237_1;
  reg                 shiftRegs_validIn_delay_238_0;
  reg                 shiftRegs_validIn_delay_238_1;
  reg                 shiftRegs_validIn_delay_239_0;
  reg                 shiftRegs_validIn_delay_239_1;
  reg                 shiftRegs_validIn_delay_240_0;
  reg                 shiftRegs_validIn_delay_240_1;
  reg                 shiftRegs_validIn_delay_241_0;
  reg                 shiftRegs_validIn_delay_241_1;
  reg                 shiftRegs_validIn_delay_242_0;
  reg                 shiftRegs_validIn_delay_242_1;
  reg                 shiftRegs_validIn_delay_243_0;
  reg                 shiftRegs_validIn_delay_243_1;
  reg                 shiftRegs_validIn_delay_244_0;
  reg                 shiftRegs_validIn_delay_244_1;
  reg                 shiftRegs_validIn_delay_245_0;
  reg                 shiftRegs_validIn_delay_245_1;
  reg                 shiftRegs_validIn_delay_246_0;
  reg                 shiftRegs_validIn_delay_246_1;
  reg                 shiftRegs_validIn_delay_247_0;
  reg                 shiftRegs_validIn_delay_247_1;
  reg                 shiftRegs_validIn_delay_248_0;
  reg                 shiftRegs_validIn_delay_248_1;
  reg                 shiftRegs_validIn_delay_249_0;
  reg                 shiftRegs_validIn_delay_249_1;
  reg                 shiftRegs_validIn_delay_250_0;
  reg                 shiftRegs_validIn_delay_250_1;
  reg                 shiftRegs_validIn_delay_251_0;
  reg                 shiftRegs_validIn_delay_251_1;
  reg                 shiftRegs_validIn_delay_252_0;
  reg                 shiftRegs_validIn_delay_252_1;
  reg                 shiftRegs_validIn_delay_253_0;
  reg                 shiftRegs_validIn_delay_253_1;
  reg                 shiftRegs_validIn_delay_254_0;
  reg                 shiftRegs_validIn_delay_254_1;
  reg                 shiftRegs_validOut_0;
  reg                 shiftRegs_validOut_1;
  reg        [15:0]   shiftRegs_addressIn_delay_1_0;
  reg        [15:0]   shiftRegs_addressIn_delay_1_1;
  reg        [15:0]   shiftRegs_addressIn_delay_2_0;
  reg        [15:0]   shiftRegs_addressIn_delay_2_1;
  reg        [15:0]   shiftRegs_addressIn_delay_3_0;
  reg        [15:0]   shiftRegs_addressIn_delay_3_1;
  reg        [15:0]   shiftRegs_addressIn_delay_4_0;
  reg        [15:0]   shiftRegs_addressIn_delay_4_1;
  reg        [15:0]   shiftRegs_addressIn_delay_5_0;
  reg        [15:0]   shiftRegs_addressIn_delay_5_1;
  reg        [15:0]   shiftRegs_addressIn_delay_6_0;
  reg        [15:0]   shiftRegs_addressIn_delay_6_1;
  reg        [15:0]   shiftRegs_addressIn_delay_7_0;
  reg        [15:0]   shiftRegs_addressIn_delay_7_1;
  reg        [15:0]   shiftRegs_addressIn_delay_8_0;
  reg        [15:0]   shiftRegs_addressIn_delay_8_1;
  reg        [15:0]   shiftRegs_addressIn_delay_9_0;
  reg        [15:0]   shiftRegs_addressIn_delay_9_1;
  reg        [15:0]   shiftRegs_addressIn_delay_10_0;
  reg        [15:0]   shiftRegs_addressIn_delay_10_1;
  reg        [15:0]   shiftRegs_addressIn_delay_11_0;
  reg        [15:0]   shiftRegs_addressIn_delay_11_1;
  reg        [15:0]   shiftRegs_addressIn_delay_12_0;
  reg        [15:0]   shiftRegs_addressIn_delay_12_1;
  reg        [15:0]   shiftRegs_addressIn_delay_13_0;
  reg        [15:0]   shiftRegs_addressIn_delay_13_1;
  reg        [15:0]   shiftRegs_addressIn_delay_14_0;
  reg        [15:0]   shiftRegs_addressIn_delay_14_1;
  reg        [15:0]   shiftRegs_addressIn_delay_15_0;
  reg        [15:0]   shiftRegs_addressIn_delay_15_1;
  reg        [15:0]   shiftRegs_addressIn_delay_16_0;
  reg        [15:0]   shiftRegs_addressIn_delay_16_1;
  reg        [15:0]   shiftRegs_addressIn_delay_17_0;
  reg        [15:0]   shiftRegs_addressIn_delay_17_1;
  reg        [15:0]   shiftRegs_addressIn_delay_18_0;
  reg        [15:0]   shiftRegs_addressIn_delay_18_1;
  reg        [15:0]   shiftRegs_addressIn_delay_19_0;
  reg        [15:0]   shiftRegs_addressIn_delay_19_1;
  reg        [15:0]   shiftRegs_addressIn_delay_20_0;
  reg        [15:0]   shiftRegs_addressIn_delay_20_1;
  reg        [15:0]   shiftRegs_addressIn_delay_21_0;
  reg        [15:0]   shiftRegs_addressIn_delay_21_1;
  reg        [15:0]   shiftRegs_addressIn_delay_22_0;
  reg        [15:0]   shiftRegs_addressIn_delay_22_1;
  reg        [15:0]   shiftRegs_addressIn_delay_23_0;
  reg        [15:0]   shiftRegs_addressIn_delay_23_1;
  reg        [15:0]   shiftRegs_addressIn_delay_24_0;
  reg        [15:0]   shiftRegs_addressIn_delay_24_1;
  reg        [15:0]   shiftRegs_addressIn_delay_25_0;
  reg        [15:0]   shiftRegs_addressIn_delay_25_1;
  reg        [15:0]   shiftRegs_addressIn_delay_26_0;
  reg        [15:0]   shiftRegs_addressIn_delay_26_1;
  reg        [15:0]   shiftRegs_addressIn_delay_27_0;
  reg        [15:0]   shiftRegs_addressIn_delay_27_1;
  reg        [15:0]   shiftRegs_addressIn_delay_28_0;
  reg        [15:0]   shiftRegs_addressIn_delay_28_1;
  reg        [15:0]   shiftRegs_addressIn_delay_29_0;
  reg        [15:0]   shiftRegs_addressIn_delay_29_1;
  reg        [15:0]   shiftRegs_addressIn_delay_30_0;
  reg        [15:0]   shiftRegs_addressIn_delay_30_1;
  reg        [15:0]   shiftRegs_addressIn_delay_31_0;
  reg        [15:0]   shiftRegs_addressIn_delay_31_1;
  reg        [15:0]   shiftRegs_addressIn_delay_32_0;
  reg        [15:0]   shiftRegs_addressIn_delay_32_1;
  reg        [15:0]   shiftRegs_addressIn_delay_33_0;
  reg        [15:0]   shiftRegs_addressIn_delay_33_1;
  reg        [15:0]   shiftRegs_addressIn_delay_34_0;
  reg        [15:0]   shiftRegs_addressIn_delay_34_1;
  reg        [15:0]   shiftRegs_addressIn_delay_35_0;
  reg        [15:0]   shiftRegs_addressIn_delay_35_1;
  reg        [15:0]   shiftRegs_addressIn_delay_36_0;
  reg        [15:0]   shiftRegs_addressIn_delay_36_1;
  reg        [15:0]   shiftRegs_addressIn_delay_37_0;
  reg        [15:0]   shiftRegs_addressIn_delay_37_1;
  reg        [15:0]   shiftRegs_addressIn_delay_38_0;
  reg        [15:0]   shiftRegs_addressIn_delay_38_1;
  reg        [15:0]   shiftRegs_addressIn_delay_39_0;
  reg        [15:0]   shiftRegs_addressIn_delay_39_1;
  reg        [15:0]   shiftRegs_addressIn_delay_40_0;
  reg        [15:0]   shiftRegs_addressIn_delay_40_1;
  reg        [15:0]   shiftRegs_addressIn_delay_41_0;
  reg        [15:0]   shiftRegs_addressIn_delay_41_1;
  reg        [15:0]   shiftRegs_addressIn_delay_42_0;
  reg        [15:0]   shiftRegs_addressIn_delay_42_1;
  reg        [15:0]   shiftRegs_addressIn_delay_43_0;
  reg        [15:0]   shiftRegs_addressIn_delay_43_1;
  reg        [15:0]   shiftRegs_addressIn_delay_44_0;
  reg        [15:0]   shiftRegs_addressIn_delay_44_1;
  reg        [15:0]   shiftRegs_addressIn_delay_45_0;
  reg        [15:0]   shiftRegs_addressIn_delay_45_1;
  reg        [15:0]   shiftRegs_addressIn_delay_46_0;
  reg        [15:0]   shiftRegs_addressIn_delay_46_1;
  reg        [15:0]   shiftRegs_addressIn_delay_47_0;
  reg        [15:0]   shiftRegs_addressIn_delay_47_1;
  reg        [15:0]   shiftRegs_addressIn_delay_48_0;
  reg        [15:0]   shiftRegs_addressIn_delay_48_1;
  reg        [15:0]   shiftRegs_addressIn_delay_49_0;
  reg        [15:0]   shiftRegs_addressIn_delay_49_1;
  reg        [15:0]   shiftRegs_addressIn_delay_50_0;
  reg        [15:0]   shiftRegs_addressIn_delay_50_1;
  reg        [15:0]   shiftRegs_addressIn_delay_51_0;
  reg        [15:0]   shiftRegs_addressIn_delay_51_1;
  reg        [15:0]   shiftRegs_addressIn_delay_52_0;
  reg        [15:0]   shiftRegs_addressIn_delay_52_1;
  reg        [15:0]   shiftRegs_addressIn_delay_53_0;
  reg        [15:0]   shiftRegs_addressIn_delay_53_1;
  reg        [15:0]   shiftRegs_addressIn_delay_54_0;
  reg        [15:0]   shiftRegs_addressIn_delay_54_1;
  reg        [15:0]   shiftRegs_addressIn_delay_55_0;
  reg        [15:0]   shiftRegs_addressIn_delay_55_1;
  reg        [15:0]   shiftRegs_addressIn_delay_56_0;
  reg        [15:0]   shiftRegs_addressIn_delay_56_1;
  reg        [15:0]   shiftRegs_addressIn_delay_57_0;
  reg        [15:0]   shiftRegs_addressIn_delay_57_1;
  reg        [15:0]   shiftRegs_addressIn_delay_58_0;
  reg        [15:0]   shiftRegs_addressIn_delay_58_1;
  reg        [15:0]   shiftRegs_addressIn_delay_59_0;
  reg        [15:0]   shiftRegs_addressIn_delay_59_1;
  reg        [15:0]   shiftRegs_addressIn_delay_60_0;
  reg        [15:0]   shiftRegs_addressIn_delay_60_1;
  reg        [15:0]   shiftRegs_addressIn_delay_61_0;
  reg        [15:0]   shiftRegs_addressIn_delay_61_1;
  reg        [15:0]   shiftRegs_addressIn_delay_62_0;
  reg        [15:0]   shiftRegs_addressIn_delay_62_1;
  reg        [15:0]   shiftRegs_addressIn_delay_63_0;
  reg        [15:0]   shiftRegs_addressIn_delay_63_1;
  reg        [15:0]   shiftRegs_addressIn_delay_64_0;
  reg        [15:0]   shiftRegs_addressIn_delay_64_1;
  reg        [15:0]   shiftRegs_addressIn_delay_65_0;
  reg        [15:0]   shiftRegs_addressIn_delay_65_1;
  reg        [15:0]   shiftRegs_addressIn_delay_66_0;
  reg        [15:0]   shiftRegs_addressIn_delay_66_1;
  reg        [15:0]   shiftRegs_addressIn_delay_67_0;
  reg        [15:0]   shiftRegs_addressIn_delay_67_1;
  reg        [15:0]   shiftRegs_addressIn_delay_68_0;
  reg        [15:0]   shiftRegs_addressIn_delay_68_1;
  reg        [15:0]   shiftRegs_addressIn_delay_69_0;
  reg        [15:0]   shiftRegs_addressIn_delay_69_1;
  reg        [15:0]   shiftRegs_addressIn_delay_70_0;
  reg        [15:0]   shiftRegs_addressIn_delay_70_1;
  reg        [15:0]   shiftRegs_addressIn_delay_71_0;
  reg        [15:0]   shiftRegs_addressIn_delay_71_1;
  reg        [15:0]   shiftRegs_addressIn_delay_72_0;
  reg        [15:0]   shiftRegs_addressIn_delay_72_1;
  reg        [15:0]   shiftRegs_addressIn_delay_73_0;
  reg        [15:0]   shiftRegs_addressIn_delay_73_1;
  reg        [15:0]   shiftRegs_addressIn_delay_74_0;
  reg        [15:0]   shiftRegs_addressIn_delay_74_1;
  reg        [15:0]   shiftRegs_addressIn_delay_75_0;
  reg        [15:0]   shiftRegs_addressIn_delay_75_1;
  reg        [15:0]   shiftRegs_addressIn_delay_76_0;
  reg        [15:0]   shiftRegs_addressIn_delay_76_1;
  reg        [15:0]   shiftRegs_addressIn_delay_77_0;
  reg        [15:0]   shiftRegs_addressIn_delay_77_1;
  reg        [15:0]   shiftRegs_addressIn_delay_78_0;
  reg        [15:0]   shiftRegs_addressIn_delay_78_1;
  reg        [15:0]   shiftRegs_addressIn_delay_79_0;
  reg        [15:0]   shiftRegs_addressIn_delay_79_1;
  reg        [15:0]   shiftRegs_addressIn_delay_80_0;
  reg        [15:0]   shiftRegs_addressIn_delay_80_1;
  reg        [15:0]   shiftRegs_addressIn_delay_81_0;
  reg        [15:0]   shiftRegs_addressIn_delay_81_1;
  reg        [15:0]   shiftRegs_addressIn_delay_82_0;
  reg        [15:0]   shiftRegs_addressIn_delay_82_1;
  reg        [15:0]   shiftRegs_addressIn_delay_83_0;
  reg        [15:0]   shiftRegs_addressIn_delay_83_1;
  reg        [15:0]   shiftRegs_addressIn_delay_84_0;
  reg        [15:0]   shiftRegs_addressIn_delay_84_1;
  reg        [15:0]   shiftRegs_addressIn_delay_85_0;
  reg        [15:0]   shiftRegs_addressIn_delay_85_1;
  reg        [15:0]   shiftRegs_addressIn_delay_86_0;
  reg        [15:0]   shiftRegs_addressIn_delay_86_1;
  reg        [15:0]   shiftRegs_addressIn_delay_87_0;
  reg        [15:0]   shiftRegs_addressIn_delay_87_1;
  reg        [15:0]   shiftRegs_addressIn_delay_88_0;
  reg        [15:0]   shiftRegs_addressIn_delay_88_1;
  reg        [15:0]   shiftRegs_addressIn_delay_89_0;
  reg        [15:0]   shiftRegs_addressIn_delay_89_1;
  reg        [15:0]   shiftRegs_addressIn_delay_90_0;
  reg        [15:0]   shiftRegs_addressIn_delay_90_1;
  reg        [15:0]   shiftRegs_addressIn_delay_91_0;
  reg        [15:0]   shiftRegs_addressIn_delay_91_1;
  reg        [15:0]   shiftRegs_addressIn_delay_92_0;
  reg        [15:0]   shiftRegs_addressIn_delay_92_1;
  reg        [15:0]   shiftRegs_addressIn_delay_93_0;
  reg        [15:0]   shiftRegs_addressIn_delay_93_1;
  reg        [15:0]   shiftRegs_addressIn_delay_94_0;
  reg        [15:0]   shiftRegs_addressIn_delay_94_1;
  reg        [15:0]   shiftRegs_addressIn_delay_95_0;
  reg        [15:0]   shiftRegs_addressIn_delay_95_1;
  reg        [15:0]   shiftRegs_addressIn_delay_96_0;
  reg        [15:0]   shiftRegs_addressIn_delay_96_1;
  reg        [15:0]   shiftRegs_addressIn_delay_97_0;
  reg        [15:0]   shiftRegs_addressIn_delay_97_1;
  reg        [15:0]   shiftRegs_addressIn_delay_98_0;
  reg        [15:0]   shiftRegs_addressIn_delay_98_1;
  reg        [15:0]   shiftRegs_addressIn_delay_99_0;
  reg        [15:0]   shiftRegs_addressIn_delay_99_1;
  reg        [15:0]   shiftRegs_addressIn_delay_100_0;
  reg        [15:0]   shiftRegs_addressIn_delay_100_1;
  reg        [15:0]   shiftRegs_addressIn_delay_101_0;
  reg        [15:0]   shiftRegs_addressIn_delay_101_1;
  reg        [15:0]   shiftRegs_addressIn_delay_102_0;
  reg        [15:0]   shiftRegs_addressIn_delay_102_1;
  reg        [15:0]   shiftRegs_addressIn_delay_103_0;
  reg        [15:0]   shiftRegs_addressIn_delay_103_1;
  reg        [15:0]   shiftRegs_addressIn_delay_104_0;
  reg        [15:0]   shiftRegs_addressIn_delay_104_1;
  reg        [15:0]   shiftRegs_addressIn_delay_105_0;
  reg        [15:0]   shiftRegs_addressIn_delay_105_1;
  reg        [15:0]   shiftRegs_addressIn_delay_106_0;
  reg        [15:0]   shiftRegs_addressIn_delay_106_1;
  reg        [15:0]   shiftRegs_addressIn_delay_107_0;
  reg        [15:0]   shiftRegs_addressIn_delay_107_1;
  reg        [15:0]   shiftRegs_addressIn_delay_108_0;
  reg        [15:0]   shiftRegs_addressIn_delay_108_1;
  reg        [15:0]   shiftRegs_addressIn_delay_109_0;
  reg        [15:0]   shiftRegs_addressIn_delay_109_1;
  reg        [15:0]   shiftRegs_addressIn_delay_110_0;
  reg        [15:0]   shiftRegs_addressIn_delay_110_1;
  reg        [15:0]   shiftRegs_addressIn_delay_111_0;
  reg        [15:0]   shiftRegs_addressIn_delay_111_1;
  reg        [15:0]   shiftRegs_addressIn_delay_112_0;
  reg        [15:0]   shiftRegs_addressIn_delay_112_1;
  reg        [15:0]   shiftRegs_addressIn_delay_113_0;
  reg        [15:0]   shiftRegs_addressIn_delay_113_1;
  reg        [15:0]   shiftRegs_addressIn_delay_114_0;
  reg        [15:0]   shiftRegs_addressIn_delay_114_1;
  reg        [15:0]   shiftRegs_addressIn_delay_115_0;
  reg        [15:0]   shiftRegs_addressIn_delay_115_1;
  reg        [15:0]   shiftRegs_addressIn_delay_116_0;
  reg        [15:0]   shiftRegs_addressIn_delay_116_1;
  reg        [15:0]   shiftRegs_addressIn_delay_117_0;
  reg        [15:0]   shiftRegs_addressIn_delay_117_1;
  reg        [15:0]   shiftRegs_addressIn_delay_118_0;
  reg        [15:0]   shiftRegs_addressIn_delay_118_1;
  reg        [15:0]   shiftRegs_addressIn_delay_119_0;
  reg        [15:0]   shiftRegs_addressIn_delay_119_1;
  reg        [15:0]   shiftRegs_addressIn_delay_120_0;
  reg        [15:0]   shiftRegs_addressIn_delay_120_1;
  reg        [15:0]   shiftRegs_addressIn_delay_121_0;
  reg        [15:0]   shiftRegs_addressIn_delay_121_1;
  reg        [15:0]   shiftRegs_addressIn_delay_122_0;
  reg        [15:0]   shiftRegs_addressIn_delay_122_1;
  reg        [15:0]   shiftRegs_addressIn_delay_123_0;
  reg        [15:0]   shiftRegs_addressIn_delay_123_1;
  reg        [15:0]   shiftRegs_addressIn_delay_124_0;
  reg        [15:0]   shiftRegs_addressIn_delay_124_1;
  reg        [15:0]   shiftRegs_addressIn_delay_125_0;
  reg        [15:0]   shiftRegs_addressIn_delay_125_1;
  reg        [15:0]   shiftRegs_addressIn_delay_126_0;
  reg        [15:0]   shiftRegs_addressIn_delay_126_1;
  reg        [15:0]   shiftRegs_addressIn_delay_127_0;
  reg        [15:0]   shiftRegs_addressIn_delay_127_1;
  reg        [15:0]   shiftRegs_addressIn_delay_128_0;
  reg        [15:0]   shiftRegs_addressIn_delay_128_1;
  reg        [15:0]   shiftRegs_addressIn_delay_129_0;
  reg        [15:0]   shiftRegs_addressIn_delay_129_1;
  reg        [15:0]   shiftRegs_addressIn_delay_130_0;
  reg        [15:0]   shiftRegs_addressIn_delay_130_1;
  reg        [15:0]   shiftRegs_addressIn_delay_131_0;
  reg        [15:0]   shiftRegs_addressIn_delay_131_1;
  reg        [15:0]   shiftRegs_addressIn_delay_132_0;
  reg        [15:0]   shiftRegs_addressIn_delay_132_1;
  reg        [15:0]   shiftRegs_addressIn_delay_133_0;
  reg        [15:0]   shiftRegs_addressIn_delay_133_1;
  reg        [15:0]   shiftRegs_addressIn_delay_134_0;
  reg        [15:0]   shiftRegs_addressIn_delay_134_1;
  reg        [15:0]   shiftRegs_addressIn_delay_135_0;
  reg        [15:0]   shiftRegs_addressIn_delay_135_1;
  reg        [15:0]   shiftRegs_addressIn_delay_136_0;
  reg        [15:0]   shiftRegs_addressIn_delay_136_1;
  reg        [15:0]   shiftRegs_addressIn_delay_137_0;
  reg        [15:0]   shiftRegs_addressIn_delay_137_1;
  reg        [15:0]   shiftRegs_addressIn_delay_138_0;
  reg        [15:0]   shiftRegs_addressIn_delay_138_1;
  reg        [15:0]   shiftRegs_addressIn_delay_139_0;
  reg        [15:0]   shiftRegs_addressIn_delay_139_1;
  reg        [15:0]   shiftRegs_addressIn_delay_140_0;
  reg        [15:0]   shiftRegs_addressIn_delay_140_1;
  reg        [15:0]   shiftRegs_addressIn_delay_141_0;
  reg        [15:0]   shiftRegs_addressIn_delay_141_1;
  reg        [15:0]   shiftRegs_addressIn_delay_142_0;
  reg        [15:0]   shiftRegs_addressIn_delay_142_1;
  reg        [15:0]   shiftRegs_addressIn_delay_143_0;
  reg        [15:0]   shiftRegs_addressIn_delay_143_1;
  reg        [15:0]   shiftRegs_addressIn_delay_144_0;
  reg        [15:0]   shiftRegs_addressIn_delay_144_1;
  reg        [15:0]   shiftRegs_addressIn_delay_145_0;
  reg        [15:0]   shiftRegs_addressIn_delay_145_1;
  reg        [15:0]   shiftRegs_addressIn_delay_146_0;
  reg        [15:0]   shiftRegs_addressIn_delay_146_1;
  reg        [15:0]   shiftRegs_addressIn_delay_147_0;
  reg        [15:0]   shiftRegs_addressIn_delay_147_1;
  reg        [15:0]   shiftRegs_addressIn_delay_148_0;
  reg        [15:0]   shiftRegs_addressIn_delay_148_1;
  reg        [15:0]   shiftRegs_addressIn_delay_149_0;
  reg        [15:0]   shiftRegs_addressIn_delay_149_1;
  reg        [15:0]   shiftRegs_addressIn_delay_150_0;
  reg        [15:0]   shiftRegs_addressIn_delay_150_1;
  reg        [15:0]   shiftRegs_addressIn_delay_151_0;
  reg        [15:0]   shiftRegs_addressIn_delay_151_1;
  reg        [15:0]   shiftRegs_addressIn_delay_152_0;
  reg        [15:0]   shiftRegs_addressIn_delay_152_1;
  reg        [15:0]   shiftRegs_addressIn_delay_153_0;
  reg        [15:0]   shiftRegs_addressIn_delay_153_1;
  reg        [15:0]   shiftRegs_addressIn_delay_154_0;
  reg        [15:0]   shiftRegs_addressIn_delay_154_1;
  reg        [15:0]   shiftRegs_addressIn_delay_155_0;
  reg        [15:0]   shiftRegs_addressIn_delay_155_1;
  reg        [15:0]   shiftRegs_addressIn_delay_156_0;
  reg        [15:0]   shiftRegs_addressIn_delay_156_1;
  reg        [15:0]   shiftRegs_addressIn_delay_157_0;
  reg        [15:0]   shiftRegs_addressIn_delay_157_1;
  reg        [15:0]   shiftRegs_addressIn_delay_158_0;
  reg        [15:0]   shiftRegs_addressIn_delay_158_1;
  reg        [15:0]   shiftRegs_addressIn_delay_159_0;
  reg        [15:0]   shiftRegs_addressIn_delay_159_1;
  reg        [15:0]   shiftRegs_addressIn_delay_160_0;
  reg        [15:0]   shiftRegs_addressIn_delay_160_1;
  reg        [15:0]   shiftRegs_addressIn_delay_161_0;
  reg        [15:0]   shiftRegs_addressIn_delay_161_1;
  reg        [15:0]   shiftRegs_addressIn_delay_162_0;
  reg        [15:0]   shiftRegs_addressIn_delay_162_1;
  reg        [15:0]   shiftRegs_addressIn_delay_163_0;
  reg        [15:0]   shiftRegs_addressIn_delay_163_1;
  reg        [15:0]   shiftRegs_addressIn_delay_164_0;
  reg        [15:0]   shiftRegs_addressIn_delay_164_1;
  reg        [15:0]   shiftRegs_addressIn_delay_165_0;
  reg        [15:0]   shiftRegs_addressIn_delay_165_1;
  reg        [15:0]   shiftRegs_addressIn_delay_166_0;
  reg        [15:0]   shiftRegs_addressIn_delay_166_1;
  reg        [15:0]   shiftRegs_addressIn_delay_167_0;
  reg        [15:0]   shiftRegs_addressIn_delay_167_1;
  reg        [15:0]   shiftRegs_addressIn_delay_168_0;
  reg        [15:0]   shiftRegs_addressIn_delay_168_1;
  reg        [15:0]   shiftRegs_addressIn_delay_169_0;
  reg        [15:0]   shiftRegs_addressIn_delay_169_1;
  reg        [15:0]   shiftRegs_addressIn_delay_170_0;
  reg        [15:0]   shiftRegs_addressIn_delay_170_1;
  reg        [15:0]   shiftRegs_addressIn_delay_171_0;
  reg        [15:0]   shiftRegs_addressIn_delay_171_1;
  reg        [15:0]   shiftRegs_addressIn_delay_172_0;
  reg        [15:0]   shiftRegs_addressIn_delay_172_1;
  reg        [15:0]   shiftRegs_addressIn_delay_173_0;
  reg        [15:0]   shiftRegs_addressIn_delay_173_1;
  reg        [15:0]   shiftRegs_addressIn_delay_174_0;
  reg        [15:0]   shiftRegs_addressIn_delay_174_1;
  reg        [15:0]   shiftRegs_addressIn_delay_175_0;
  reg        [15:0]   shiftRegs_addressIn_delay_175_1;
  reg        [15:0]   shiftRegs_addressIn_delay_176_0;
  reg        [15:0]   shiftRegs_addressIn_delay_176_1;
  reg        [15:0]   shiftRegs_addressIn_delay_177_0;
  reg        [15:0]   shiftRegs_addressIn_delay_177_1;
  reg        [15:0]   shiftRegs_addressIn_delay_178_0;
  reg        [15:0]   shiftRegs_addressIn_delay_178_1;
  reg        [15:0]   shiftRegs_addressIn_delay_179_0;
  reg        [15:0]   shiftRegs_addressIn_delay_179_1;
  reg        [15:0]   shiftRegs_addressIn_delay_180_0;
  reg        [15:0]   shiftRegs_addressIn_delay_180_1;
  reg        [15:0]   shiftRegs_addressIn_delay_181_0;
  reg        [15:0]   shiftRegs_addressIn_delay_181_1;
  reg        [15:0]   shiftRegs_addressIn_delay_182_0;
  reg        [15:0]   shiftRegs_addressIn_delay_182_1;
  reg        [15:0]   shiftRegs_addressIn_delay_183_0;
  reg        [15:0]   shiftRegs_addressIn_delay_183_1;
  reg        [15:0]   shiftRegs_addressIn_delay_184_0;
  reg        [15:0]   shiftRegs_addressIn_delay_184_1;
  reg        [15:0]   shiftRegs_addressIn_delay_185_0;
  reg        [15:0]   shiftRegs_addressIn_delay_185_1;
  reg        [15:0]   shiftRegs_addressIn_delay_186_0;
  reg        [15:0]   shiftRegs_addressIn_delay_186_1;
  reg        [15:0]   shiftRegs_addressIn_delay_187_0;
  reg        [15:0]   shiftRegs_addressIn_delay_187_1;
  reg        [15:0]   shiftRegs_addressIn_delay_188_0;
  reg        [15:0]   shiftRegs_addressIn_delay_188_1;
  reg        [15:0]   shiftRegs_addressIn_delay_189_0;
  reg        [15:0]   shiftRegs_addressIn_delay_189_1;
  reg        [15:0]   shiftRegs_addressIn_delay_190_0;
  reg        [15:0]   shiftRegs_addressIn_delay_190_1;
  reg        [15:0]   shiftRegs_addressIn_delay_191_0;
  reg        [15:0]   shiftRegs_addressIn_delay_191_1;
  reg        [15:0]   shiftRegs_addressIn_delay_192_0;
  reg        [15:0]   shiftRegs_addressIn_delay_192_1;
  reg        [15:0]   shiftRegs_addressIn_delay_193_0;
  reg        [15:0]   shiftRegs_addressIn_delay_193_1;
  reg        [15:0]   shiftRegs_addressIn_delay_194_0;
  reg        [15:0]   shiftRegs_addressIn_delay_194_1;
  reg        [15:0]   shiftRegs_addressIn_delay_195_0;
  reg        [15:0]   shiftRegs_addressIn_delay_195_1;
  reg        [15:0]   shiftRegs_addressIn_delay_196_0;
  reg        [15:0]   shiftRegs_addressIn_delay_196_1;
  reg        [15:0]   shiftRegs_addressIn_delay_197_0;
  reg        [15:0]   shiftRegs_addressIn_delay_197_1;
  reg        [15:0]   shiftRegs_addressIn_delay_198_0;
  reg        [15:0]   shiftRegs_addressIn_delay_198_1;
  reg        [15:0]   shiftRegs_addressIn_delay_199_0;
  reg        [15:0]   shiftRegs_addressIn_delay_199_1;
  reg        [15:0]   shiftRegs_addressIn_delay_200_0;
  reg        [15:0]   shiftRegs_addressIn_delay_200_1;
  reg        [15:0]   shiftRegs_addressIn_delay_201_0;
  reg        [15:0]   shiftRegs_addressIn_delay_201_1;
  reg        [15:0]   shiftRegs_addressIn_delay_202_0;
  reg        [15:0]   shiftRegs_addressIn_delay_202_1;
  reg        [15:0]   shiftRegs_addressIn_delay_203_0;
  reg        [15:0]   shiftRegs_addressIn_delay_203_1;
  reg        [15:0]   shiftRegs_addressIn_delay_204_0;
  reg        [15:0]   shiftRegs_addressIn_delay_204_1;
  reg        [15:0]   shiftRegs_addressIn_delay_205_0;
  reg        [15:0]   shiftRegs_addressIn_delay_205_1;
  reg        [15:0]   shiftRegs_addressIn_delay_206_0;
  reg        [15:0]   shiftRegs_addressIn_delay_206_1;
  reg        [15:0]   shiftRegs_addressIn_delay_207_0;
  reg        [15:0]   shiftRegs_addressIn_delay_207_1;
  reg        [15:0]   shiftRegs_addressIn_delay_208_0;
  reg        [15:0]   shiftRegs_addressIn_delay_208_1;
  reg        [15:0]   shiftRegs_addressIn_delay_209_0;
  reg        [15:0]   shiftRegs_addressIn_delay_209_1;
  reg        [15:0]   shiftRegs_addressIn_delay_210_0;
  reg        [15:0]   shiftRegs_addressIn_delay_210_1;
  reg        [15:0]   shiftRegs_addressIn_delay_211_0;
  reg        [15:0]   shiftRegs_addressIn_delay_211_1;
  reg        [15:0]   shiftRegs_addressIn_delay_212_0;
  reg        [15:0]   shiftRegs_addressIn_delay_212_1;
  reg        [15:0]   shiftRegs_addressIn_delay_213_0;
  reg        [15:0]   shiftRegs_addressIn_delay_213_1;
  reg        [15:0]   shiftRegs_addressIn_delay_214_0;
  reg        [15:0]   shiftRegs_addressIn_delay_214_1;
  reg        [15:0]   shiftRegs_addressIn_delay_215_0;
  reg        [15:0]   shiftRegs_addressIn_delay_215_1;
  reg        [15:0]   shiftRegs_addressIn_delay_216_0;
  reg        [15:0]   shiftRegs_addressIn_delay_216_1;
  reg        [15:0]   shiftRegs_addressIn_delay_217_0;
  reg        [15:0]   shiftRegs_addressIn_delay_217_1;
  reg        [15:0]   shiftRegs_addressIn_delay_218_0;
  reg        [15:0]   shiftRegs_addressIn_delay_218_1;
  reg        [15:0]   shiftRegs_addressIn_delay_219_0;
  reg        [15:0]   shiftRegs_addressIn_delay_219_1;
  reg        [15:0]   shiftRegs_addressIn_delay_220_0;
  reg        [15:0]   shiftRegs_addressIn_delay_220_1;
  reg        [15:0]   shiftRegs_addressIn_delay_221_0;
  reg        [15:0]   shiftRegs_addressIn_delay_221_1;
  reg        [15:0]   shiftRegs_addressIn_delay_222_0;
  reg        [15:0]   shiftRegs_addressIn_delay_222_1;
  reg        [15:0]   shiftRegs_addressIn_delay_223_0;
  reg        [15:0]   shiftRegs_addressIn_delay_223_1;
  reg        [15:0]   shiftRegs_addressIn_delay_224_0;
  reg        [15:0]   shiftRegs_addressIn_delay_224_1;
  reg        [15:0]   shiftRegs_addressIn_delay_225_0;
  reg        [15:0]   shiftRegs_addressIn_delay_225_1;
  reg        [15:0]   shiftRegs_addressIn_delay_226_0;
  reg        [15:0]   shiftRegs_addressIn_delay_226_1;
  reg        [15:0]   shiftRegs_addressIn_delay_227_0;
  reg        [15:0]   shiftRegs_addressIn_delay_227_1;
  reg        [15:0]   shiftRegs_addressIn_delay_228_0;
  reg        [15:0]   shiftRegs_addressIn_delay_228_1;
  reg        [15:0]   shiftRegs_addressIn_delay_229_0;
  reg        [15:0]   shiftRegs_addressIn_delay_229_1;
  reg        [15:0]   shiftRegs_addressIn_delay_230_0;
  reg        [15:0]   shiftRegs_addressIn_delay_230_1;
  reg        [15:0]   shiftRegs_addressIn_delay_231_0;
  reg        [15:0]   shiftRegs_addressIn_delay_231_1;
  reg        [15:0]   shiftRegs_addressIn_delay_232_0;
  reg        [15:0]   shiftRegs_addressIn_delay_232_1;
  reg        [15:0]   shiftRegs_addressIn_delay_233_0;
  reg        [15:0]   shiftRegs_addressIn_delay_233_1;
  reg        [15:0]   shiftRegs_addressIn_delay_234_0;
  reg        [15:0]   shiftRegs_addressIn_delay_234_1;
  reg        [15:0]   shiftRegs_addressIn_delay_235_0;
  reg        [15:0]   shiftRegs_addressIn_delay_235_1;
  reg        [15:0]   shiftRegs_addressIn_delay_236_0;
  reg        [15:0]   shiftRegs_addressIn_delay_236_1;
  reg        [15:0]   shiftRegs_addressIn_delay_237_0;
  reg        [15:0]   shiftRegs_addressIn_delay_237_1;
  reg        [15:0]   shiftRegs_addressIn_delay_238_0;
  reg        [15:0]   shiftRegs_addressIn_delay_238_1;
  reg        [15:0]   shiftRegs_addressIn_delay_239_0;
  reg        [15:0]   shiftRegs_addressIn_delay_239_1;
  reg        [15:0]   shiftRegs_addressIn_delay_240_0;
  reg        [15:0]   shiftRegs_addressIn_delay_240_1;
  reg        [15:0]   shiftRegs_addressIn_delay_241_0;
  reg        [15:0]   shiftRegs_addressIn_delay_241_1;
  reg        [15:0]   shiftRegs_addressIn_delay_242_0;
  reg        [15:0]   shiftRegs_addressIn_delay_242_1;
  reg        [15:0]   shiftRegs_addressIn_delay_243_0;
  reg        [15:0]   shiftRegs_addressIn_delay_243_1;
  reg        [15:0]   shiftRegs_addressIn_delay_244_0;
  reg        [15:0]   shiftRegs_addressIn_delay_244_1;
  reg        [15:0]   shiftRegs_addressIn_delay_245_0;
  reg        [15:0]   shiftRegs_addressIn_delay_245_1;
  reg        [15:0]   shiftRegs_addressIn_delay_246_0;
  reg        [15:0]   shiftRegs_addressIn_delay_246_1;
  reg        [15:0]   shiftRegs_addressIn_delay_247_0;
  reg        [15:0]   shiftRegs_addressIn_delay_247_1;
  reg        [15:0]   shiftRegs_addressIn_delay_248_0;
  reg        [15:0]   shiftRegs_addressIn_delay_248_1;
  reg        [15:0]   shiftRegs_addressIn_delay_249_0;
  reg        [15:0]   shiftRegs_addressIn_delay_249_1;
  reg        [15:0]   shiftRegs_addressIn_delay_250_0;
  reg        [15:0]   shiftRegs_addressIn_delay_250_1;
  reg        [15:0]   shiftRegs_addressIn_delay_251_0;
  reg        [15:0]   shiftRegs_addressIn_delay_251_1;
  reg        [15:0]   shiftRegs_addressIn_delay_252_0;
  reg        [15:0]   shiftRegs_addressIn_delay_252_1;
  reg        [15:0]   shiftRegs_addressIn_delay_253_0;
  reg        [15:0]   shiftRegs_addressIn_delay_253_1;
  reg        [15:0]   shiftRegs_addressIn_delay_254_0;
  reg        [15:0]   shiftRegs_addressIn_delay_254_1;
  reg        [15:0]   shiftRegs_addressOut_0;
  reg        [15:0]   shiftRegs_addressOut_1;
  reg                 shiftRegs_validOut_delay_1_0;
  reg                 shiftRegs_validOut_delay_1_1;
  reg                 shiftRegs_validOut_delay_2_0;
  reg                 shiftRegs_validOut_delay_2_1;
  reg                 shiftRegs_validOut_delay_3_0;
  reg                 shiftRegs_validOut_delay_3_1;
  reg                 shiftRegs_validOut_delay_4_0;
  reg                 shiftRegs_validOut_delay_4_1;
  reg                 shiftRegs_validOutFull_0;
  reg                 shiftRegs_validOutFull_1;
  reg        [15:0]   shiftRegs_addressOut_delay_1_0;
  reg        [15:0]   shiftRegs_addressOut_delay_1_1;
  reg        [15:0]   shiftRegs_addressOut_delay_2_0;
  reg        [15:0]   shiftRegs_addressOut_delay_2_1;
  reg        [15:0]   shiftRegs_addressOut_delay_3_0;
  reg        [15:0]   shiftRegs_addressOut_delay_3_1;
  reg        [15:0]   shiftRegs_addressOut_delay_4_0;
  reg        [15:0]   shiftRegs_addressOut_delay_4_1;
  reg        [15:0]   shiftRegs_addressOutFull_0;
  reg        [15:0]   shiftRegs_addressOutFull_1;
  reg                 outputValid;
  reg        [376:0]  pAddPort_0_s_regNext_X;
  reg        [376:0]  pAddPort_0_s_regNext_Y;
  reg        [376:0]  pAddPort_0_s_regNext_Z;
  reg        [376:0]  pAddPort_0_s_regNext_T;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg                 flushing_flushCnt_willIncrement;
  wire                flushing_flushCnt_willClear;
  reg        [15:0]   flushing_flushCnt_valueNext;
  reg        [15:0]   flushing_flushCnt_value;
  reg                 flushing_flushCnt_willOverflowIfInc;
  wire                flushing_flushCnt_willOverflow;
  reg                 stage1_NCnt_willIncrement;
  reg                 stage1_NCnt_willClear;
  reg        [31:0]   stage1_NCnt_valueNext;
  reg        [31:0]   stage1_NCnt_value;
  reg                 stage1_NCnt_willOverflowIfInc;
  wire                stage1_NCnt_willOverflow;
  reg                 stage1_GCnt_willIncrement;
  wire                stage1_GCnt_willClear;
  reg        [3:0]    stage1_GCnt_valueNext;
  reg        [3:0]    stage1_GCnt_value;
  reg                 stage1_GCnt_willOverflowIfInc;
  wire                stage1_GCnt_willOverflow;
  reg                 stage1_waitReg;
  reg                 stage1_emptyCnt_willIncrement;
  reg                 stage1_emptyCnt_willClear;
  reg        [8:0]    stage1_emptyCnt_valueNext;
  reg        [8:0]    stage1_emptyCnt_value;
  reg                 stage1_emptyCnt_willOverflowIfInc;
  wire                stage1_emptyCnt_willOverflow;
  reg                 stage1_needAdd1_0;
  wire       [25:0]   _zz_stage1_inputBarrelID_0;
  wire       [13:0]   stage1_inputBarrelID_0;
  wire       [13:0]   stage1_inputBarrelID_1;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0;
  wire       [11:0]   stage1_inputBarrelIDAbs_0;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_1;
  wire       [11:0]   stage1_inputBarrelIDAbs_1;
  reg                 _zz_stage1_inputValid_0;
  reg                 _zz_stage1_inputValid_0_1;
  reg                 _zz_stage1_inputValid_0_2;
  reg                 _zz_stage1_inputValid_0_3;
  reg                 _zz_stage1_inputValid_0_4;
  reg                 stage1_inputValid_0;
  reg                 _zz_stage1_inputValid_1;
  reg                 _zz_stage1_inputValid_1_1;
  reg                 _zz_stage1_inputValid_1_2;
  reg                 _zz_stage1_inputValid_1_3;
  reg                 _zz_stage1_inputValid_1_4;
  reg                 stage1_inputValid_1;
  reg        [15:0]   _zz_stage1_inputAddress_0;
  reg        [15:0]   _zz_stage1_inputAddress_0_1;
  reg        [15:0]   _zz_stage1_inputAddress_0_2;
  reg        [15:0]   _zz_stage1_inputAddress_0_3;
  reg        [15:0]   _zz_stage1_inputAddress_0_4;
  reg        [15:0]   stage1_inputAddress_0;
  reg        [15:0]   _zz_stage1_inputAddress_1;
  reg        [15:0]   _zz_stage1_inputAddress_1_1;
  reg        [15:0]   _zz_stage1_inputAddress_1_2;
  reg        [15:0]   _zz_stage1_inputAddress_1_3;
  reg        [15:0]   _zz_stage1_inputAddress_1_4;
  reg        [15:0]   stage1_inputAddress_1;
  reg                 _zz_stage1_inputData_0_X;
  reg                 _zz_stage1_inputData_0_X_1;
  reg                 _zz_stage1_inputData_0_X_2;
  reg                 _zz_stage1_inputData_0_X_3;
  reg                 _zz_stage1_inputData_0_X_4;
  reg                 _zz_stage1_inputData_0_X_5;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_T;
  wire       [376:0]  stage1_inputData_0_X;
  wire       [376:0]  stage1_inputData_0_Y;
  wire       [376:0]  stage1_inputData_0_Z;
  wire       [376:0]  stage1_inputData_0_T;
  reg                 _zz_stage1_inputData_1_X;
  reg                 _zz_stage1_inputData_1_X_1;
  reg                 _zz_stage1_inputData_1_X_2;
  reg                 _zz_stage1_inputData_1_X_3;
  reg                 _zz_stage1_inputData_1_X_4;
  reg                 _zz_stage1_inputData_1_X_5;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_X_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_T_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_X_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_T_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_X_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_T_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_X_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_T_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_X_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_T_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_X_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z_1;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_T_1;
  wire       [376:0]  stage1_inputData_1_X;
  wire       [376:0]  stage1_inputData_1_Y;
  wire       [376:0]  stage1_inputData_1_Z;
  wire       [376:0]  stage1_inputData_1_T;
  reg                 stage2_wCnt_willDecrement;
  wire                stage2_wCnt_willClear;
  reg        [11:0]   stage2_wCnt_valueNext;
  reg        [11:0]   stage2_wCnt_value;
  reg                 stage2_wCnt_willUnderflowIfDec;
  wire                stage2_wCnt_willUnderflow;
  reg                 stage2_GCnt_willIncrement;
  wire                stage2_GCnt_willClear;
  reg        [3:0]    stage2_GCnt_valueNext;
  reg        [3:0]    stage2_GCnt_value;
  reg                 stage2_GCnt_willOverflowIfInc;
  wire                stage2_GCnt_willOverflow;
  reg                 stage2_calCnt_willDecrement;
  wire                stage2_calCnt_willClear;
  reg        [1:0]    stage2_calCnt_valueNext;
  reg        [1:0]    stage2_calCnt_value;
  reg                 stage2_calCnt_willUnderflowIfDec;
  wire                stage2_calCnt_willUnderflow;
  reg                 stage2_waitReg;
  reg                 stage2_waitCnt_willIncrement;
  wire                stage2_waitCnt_willClear;
  reg        [8:0]    stage2_waitCnt_valueNext;
  reg        [8:0]    stage2_waitCnt_value;
  reg                 stage2_waitCnt_willOverflowIfInc;
  wire                stage2_waitCnt_willOverflow;
  reg                 stage3_GCnt_willDecrement;
  wire                stage3_GCnt_willClear;
  reg        [3:0]    stage3_GCnt_valueNext;
  reg        [3:0]    stage3_GCnt_value;
  reg                 stage3_GCnt_willUnderflowIfDec;
  wire                stage3_GCnt_willUnderflow;
  reg                 stage3_doubleCnt_willIncrement;
  wire                stage3_doubleCnt_willClear;
  reg        [4:0]    stage3_doubleCnt_valueNext;
  reg        [4:0]    stage3_doubleCnt_value;
  reg                 stage3_doubleCnt_willOverflowIfInc;
  wire                stage3_doubleCnt_willOverflow;
  reg                 stage3_doubleWaitCnt_willIncrement;
  wire                stage3_doubleWaitCnt_willClear;
  reg        [8:0]    stage3_doubleWaitCnt_valueNext;
  reg        [8:0]    stage3_doubleWaitCnt_value;
  reg                 stage3_doubleWaitCnt_willOverflowIfInc;
  wire                stage3_doubleWaitCnt_willOverflow;
  reg                 stage3_addReg;
  reg                 stage3_addWaitCnt_willIncrement;
  wire                stage3_addWaitCnt_willClear;
  reg        [8:0]    stage3_addWaitCnt_valueNext;
  reg        [8:0]    stage3_addWaitCnt_value;
  reg                 stage3_addWaitCnt_willOverflowIfInc;
  wire                stage3_addWaitCnt_willOverflow;
  reg                 stage3Final_doubleCnt_willIncrement;
  wire                stage3Final_doubleCnt_willClear;
  reg        [3:0]    stage3Final_doubleCnt_valueNext;
  reg        [3:0]    stage3Final_doubleCnt_value;
  reg                 stage3Final_doubleCnt_willOverflowIfInc;
  wire                stage3Final_doubleCnt_willOverflow;
  reg                 stage3Final_doubleWaitCnt_willIncrement;
  wire                stage3Final_doubleWaitCnt_willClear;
  reg        [8:0]    stage3Final_doubleWaitCnt_valueNext;
  reg        [8:0]    stage3Final_doubleWaitCnt_value;
  reg                 stage3Final_doubleWaitCnt_willOverflowIfInc;
  wire                stage3Final_doubleWaitCnt_willOverflow;
  reg                 stage3Final_addReg;
  reg                 stage3Final_addWaitCnt_willIncrement;
  wire                stage3Final_addWaitCnt_willClear;
  reg        [8:0]    stage3Final_addWaitCnt_valueNext;
  reg        [8:0]    stage3Final_addWaitCnt_value;
  reg                 stage3Final_addWaitCnt_willOverflowIfInc;
  wire                stage3Final_addWaitCnt_willOverflow;
  reg        [0:0]    stage3Final_pAddShr;
  reg        [4:0]    fsm_stateReg;
  reg        [4:0]    fsm_stateNext;
  reg                 stage1_inputValid_0_delay_1;
  reg                 stage1_inputValid_0_delay_2;
  reg                 stage1_inputValid_0_delay_3;
  reg                 stage1_inputValid_0_delay_4;
  reg                 stage1_inputValid_0_delay_5;
  reg        [15:0]   stage1_inputAddress_0_delay_1;
  reg        [15:0]   stage1_inputAddress_0_delay_2;
  reg        [15:0]   stage1_inputAddress_0_delay_3;
  reg        [15:0]   stage1_inputAddress_0_delay_4;
  reg        [15:0]   stage1_inputAddress_0_delay_5;
  reg        [376:0]  stage1_inputData_0_delay_1_X;
  reg        [376:0]  stage1_inputData_0_delay_1_Y;
  reg        [376:0]  stage1_inputData_0_delay_1_Z;
  reg        [376:0]  stage1_inputData_0_delay_1_T;
  reg        [376:0]  stage1_inputData_0_delay_2_X;
  reg        [376:0]  stage1_inputData_0_delay_2_Y;
  reg        [376:0]  stage1_inputData_0_delay_2_Z;
  reg        [376:0]  stage1_inputData_0_delay_2_T;
  reg        [376:0]  stage1_inputData_0_delay_3_X;
  reg        [376:0]  stage1_inputData_0_delay_3_Y;
  reg        [376:0]  stage1_inputData_0_delay_3_Z;
  reg        [376:0]  stage1_inputData_0_delay_3_T;
  reg        [376:0]  stage1_inputData_0_delay_4_X;
  reg        [376:0]  stage1_inputData_0_delay_4_Y;
  reg        [376:0]  stage1_inputData_0_delay_4_Z;
  reg        [376:0]  stage1_inputData_0_delay_4_T;
  reg        [376:0]  stage1_inputData_0_delay_5_X;
  reg        [376:0]  stage1_inputData_0_delay_5_Y;
  reg        [376:0]  stage1_inputData_0_delay_5_Z;
  reg        [376:0]  stage1_inputData_0_delay_5_T;
  reg                 _zz_io_dataIn_0_valid;
  reg                 _zz_io_dataIn_0_valid_1;
  reg                 _zz_io_dataIn_0_valid_2;
  reg                 _zz_io_dataIn_0_valid_3;
  reg                 _zz_io_dataIn_0_valid_4;
  reg                 _zz_io_dataIn_0_valid_5;
  reg                 _zz_io_dataIn_0_valid_6;
  reg                 _zz_io_dataIn_0_valid_7;
  reg                 _zz_io_dataIn_0_valid_8;
  reg                 _zz_io_dataIn_0_valid_9;
  reg                 _zz_io_dataIn_0_valid_10;
  reg                 _zz_io_dataIn_0_valid_11;
  reg                 _zz_io_dataIn_0_valid_12;
  reg                 _zz_io_dataIn_0_valid_13;
  reg                 _zz_io_dataIn_0_valid_14;
  reg                 _zz_io_dataIn_0_valid_15;
  reg                 _zz_io_dataIn_0_valid_16;
  reg                 _zz_io_dataIn_0_valid_17;
  reg                 _zz_io_dataIn_0_valid_18;
  reg                 _zz_io_dataIn_0_valid_19;
  reg                 _zz_io_dataIn_0_valid_20;
  reg                 _zz_io_dataIn_0_valid_21;
  reg                 _zz_io_dataIn_0_valid_22;
  reg                 _zz_io_dataIn_0_valid_23;
  reg                 _zz_io_dataIn_0_valid_24;
  reg                 _zz_io_dataIn_0_valid_25;
  reg                 _zz_io_dataIn_0_valid_26;
  reg                 _zz_io_dataIn_0_valid_27;
  reg                 _zz_io_dataIn_0_valid_28;
  reg                 _zz_io_dataIn_0_valid_29;
  reg                 _zz_io_dataIn_0_valid_30;
  reg                 _zz_io_dataIn_0_valid_31;
  reg                 _zz_io_dataIn_0_valid_32;
  reg                 _zz_io_dataIn_0_valid_33;
  reg                 _zz_io_dataIn_0_valid_34;
  reg                 _zz_io_dataIn_0_payload_a_X;
  reg                 _zz_io_dataIn_0_payload_a_X_1;
  reg                 _zz_io_dataIn_0_payload_a_X_2;
  reg                 _zz_io_dataIn_0_payload_a_X_3;
  reg                 _zz_io_dataIn_0_payload_a_X_4;
  reg                 _zz_io_dataIn_0_payload_a_X_5;
  reg                 _zz_io_dataIn_0_payload_a_X_6;
  reg                 _zz_io_dataIn_0_payload_a_X_7;
  reg                 _zz_io_dataIn_0_payload_a_X_8;
  reg                 _zz_io_dataIn_0_payload_a_X_9;
  reg                 _zz_io_dataIn_0_payload_a_X_10;
  reg                 _zz_io_dataIn_0_payload_a_X_11;
  reg                 _zz_io_dataIn_0_payload_a_X_12;
  reg                 _zz_io_dataIn_0_payload_a_X_13;
  reg                 _zz_io_dataIn_0_payload_a_X_14;
  reg                 _zz_io_dataIn_0_payload_a_X_15;
  reg                 _zz_io_dataIn_0_payload_a_X_16;
  reg                 _zz_io_dataIn_0_payload_a_X_17;
  reg                 _zz_io_dataIn_0_payload_a_X_18;
  reg                 _zz_io_dataIn_0_payload_a_X_19;
  reg                 _zz_io_dataIn_0_payload_a_X_20;
  reg                 _zz_io_dataIn_0_payload_a_X_21;
  reg                 _zz_io_dataIn_0_payload_a_X_22;
  reg                 _zz_io_dataIn_0_payload_a_X_23;
  reg                 _zz_io_dataIn_0_payload_a_X_24;
  reg                 _zz_io_dataIn_0_payload_a_X_25;
  reg                 _zz_io_dataIn_0_payload_a_X_26;
  reg                 _zz_io_dataIn_0_payload_a_X_27;
  reg                 _zz_io_dataIn_0_payload_a_X_28;
  reg                 _zz_io_dataIn_0_payload_a_X_29;
  reg                 _zz_io_dataIn_0_payload_a_X_30;
  reg                 _zz_io_dataIn_0_payload_a_X_31;
  reg                 _zz_io_dataIn_0_payload_a_X_32;
  reg                 _zz_io_dataIn_0_payload_a_X_33;
  reg                 _zz_io_dataIn_0_payload_a_X_34;
  reg        [376:0]  stage1_inputData_0_delay_1_X_1;
  reg        [376:0]  stage1_inputData_0_delay_1_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_1_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_1_T_1;
  reg        [376:0]  stage1_inputData_0_delay_2_X_1;
  reg        [376:0]  stage1_inputData_0_delay_2_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_2_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_2_T_1;
  reg        [376:0]  stage1_inputData_0_delay_3_X_1;
  reg        [376:0]  stage1_inputData_0_delay_3_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_3_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_3_T_1;
  reg        [376:0]  stage1_inputData_0_delay_4_X_1;
  reg        [376:0]  stage1_inputData_0_delay_4_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_4_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_4_T_1;
  reg        [376:0]  stage1_inputData_0_delay_5_X_1;
  reg        [376:0]  stage1_inputData_0_delay_5_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_5_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_5_T_1;
  reg        [376:0]  stage1_inputData_0_delay_6_X;
  reg        [376:0]  stage1_inputData_0_delay_6_Y;
  reg        [376:0]  stage1_inputData_0_delay_6_Z;
  reg        [376:0]  stage1_inputData_0_delay_6_T;
  reg        [376:0]  stage1_inputData_0_delay_7_X;
  reg        [376:0]  stage1_inputData_0_delay_7_Y;
  reg        [376:0]  stage1_inputData_0_delay_7_Z;
  reg        [376:0]  stage1_inputData_0_delay_7_T;
  reg        [376:0]  stage1_inputData_0_delay_8_X;
  reg        [376:0]  stage1_inputData_0_delay_8_Y;
  reg        [376:0]  stage1_inputData_0_delay_8_Z;
  reg        [376:0]  stage1_inputData_0_delay_8_T;
  reg        [376:0]  stage1_inputData_0_delay_9_X;
  reg        [376:0]  stage1_inputData_0_delay_9_Y;
  reg        [376:0]  stage1_inputData_0_delay_9_Z;
  reg        [376:0]  stage1_inputData_0_delay_9_T;
  reg        [376:0]  stage1_inputData_0_delay_10_X;
  reg        [376:0]  stage1_inputData_0_delay_10_Y;
  reg        [376:0]  stage1_inputData_0_delay_10_Z;
  reg        [376:0]  stage1_inputData_0_delay_10_T;
  reg        [376:0]  stage1_inputData_0_delay_11_X;
  reg        [376:0]  stage1_inputData_0_delay_11_Y;
  reg        [376:0]  stage1_inputData_0_delay_11_Z;
  reg        [376:0]  stage1_inputData_0_delay_11_T;
  reg        [376:0]  stage1_inputData_0_delay_12_X;
  reg        [376:0]  stage1_inputData_0_delay_12_Y;
  reg        [376:0]  stage1_inputData_0_delay_12_Z;
  reg        [376:0]  stage1_inputData_0_delay_12_T;
  reg        [376:0]  stage1_inputData_0_delay_13_X;
  reg        [376:0]  stage1_inputData_0_delay_13_Y;
  reg        [376:0]  stage1_inputData_0_delay_13_Z;
  reg        [376:0]  stage1_inputData_0_delay_13_T;
  reg        [376:0]  stage1_inputData_0_delay_14_X;
  reg        [376:0]  stage1_inputData_0_delay_14_Y;
  reg        [376:0]  stage1_inputData_0_delay_14_Z;
  reg        [376:0]  stage1_inputData_0_delay_14_T;
  reg        [376:0]  stage1_inputData_0_delay_15_X;
  reg        [376:0]  stage1_inputData_0_delay_15_Y;
  reg        [376:0]  stage1_inputData_0_delay_15_Z;
  reg        [376:0]  stage1_inputData_0_delay_15_T;
  reg        [376:0]  stage1_inputData_0_delay_16_X;
  reg        [376:0]  stage1_inputData_0_delay_16_Y;
  reg        [376:0]  stage1_inputData_0_delay_16_Z;
  reg        [376:0]  stage1_inputData_0_delay_16_T;
  reg        [376:0]  stage1_inputData_0_delay_17_X;
  reg        [376:0]  stage1_inputData_0_delay_17_Y;
  reg        [376:0]  stage1_inputData_0_delay_17_Z;
  reg        [376:0]  stage1_inputData_0_delay_17_T;
  reg        [376:0]  stage1_inputData_0_delay_18_X;
  reg        [376:0]  stage1_inputData_0_delay_18_Y;
  reg        [376:0]  stage1_inputData_0_delay_18_Z;
  reg        [376:0]  stage1_inputData_0_delay_18_T;
  reg        [376:0]  stage1_inputData_0_delay_19_X;
  reg        [376:0]  stage1_inputData_0_delay_19_Y;
  reg        [376:0]  stage1_inputData_0_delay_19_Z;
  reg        [376:0]  stage1_inputData_0_delay_19_T;
  reg        [376:0]  stage1_inputData_0_delay_20_X;
  reg        [376:0]  stage1_inputData_0_delay_20_Y;
  reg        [376:0]  stage1_inputData_0_delay_20_Z;
  reg        [376:0]  stage1_inputData_0_delay_20_T;
  reg        [376:0]  stage1_inputData_0_delay_21_X;
  reg        [376:0]  stage1_inputData_0_delay_21_Y;
  reg        [376:0]  stage1_inputData_0_delay_21_Z;
  reg        [376:0]  stage1_inputData_0_delay_21_T;
  reg        [376:0]  stage1_inputData_0_delay_22_X;
  reg        [376:0]  stage1_inputData_0_delay_22_Y;
  reg        [376:0]  stage1_inputData_0_delay_22_Z;
  reg        [376:0]  stage1_inputData_0_delay_22_T;
  reg        [376:0]  stage1_inputData_0_delay_23_X;
  reg        [376:0]  stage1_inputData_0_delay_23_Y;
  reg        [376:0]  stage1_inputData_0_delay_23_Z;
  reg        [376:0]  stage1_inputData_0_delay_23_T;
  reg        [376:0]  stage1_inputData_0_delay_24_X;
  reg        [376:0]  stage1_inputData_0_delay_24_Y;
  reg        [376:0]  stage1_inputData_0_delay_24_Z;
  reg        [376:0]  stage1_inputData_0_delay_24_T;
  reg        [376:0]  stage1_inputData_0_delay_25_X;
  reg        [376:0]  stage1_inputData_0_delay_25_Y;
  reg        [376:0]  stage1_inputData_0_delay_25_Z;
  reg        [376:0]  stage1_inputData_0_delay_25_T;
  reg        [376:0]  stage1_inputData_0_delay_26_X;
  reg        [376:0]  stage1_inputData_0_delay_26_Y;
  reg        [376:0]  stage1_inputData_0_delay_26_Z;
  reg        [376:0]  stage1_inputData_0_delay_26_T;
  reg        [376:0]  stage1_inputData_0_delay_27_X;
  reg        [376:0]  stage1_inputData_0_delay_27_Y;
  reg        [376:0]  stage1_inputData_0_delay_27_Z;
  reg        [376:0]  stage1_inputData_0_delay_27_T;
  reg        [376:0]  stage1_inputData_0_delay_28_X;
  reg        [376:0]  stage1_inputData_0_delay_28_Y;
  reg        [376:0]  stage1_inputData_0_delay_28_Z;
  reg        [376:0]  stage1_inputData_0_delay_28_T;
  reg        [376:0]  stage1_inputData_0_delay_29_X;
  reg        [376:0]  stage1_inputData_0_delay_29_Y;
  reg        [376:0]  stage1_inputData_0_delay_29_Z;
  reg        [376:0]  stage1_inputData_0_delay_29_T;
  reg        [376:0]  stage1_inputData_0_delay_30_X;
  reg        [376:0]  stage1_inputData_0_delay_30_Y;
  reg        [376:0]  stage1_inputData_0_delay_30_Z;
  reg        [376:0]  stage1_inputData_0_delay_30_T;
  reg        [376:0]  stage1_inputData_0_delay_31_X;
  reg        [376:0]  stage1_inputData_0_delay_31_Y;
  reg        [376:0]  stage1_inputData_0_delay_31_Z;
  reg        [376:0]  stage1_inputData_0_delay_31_T;
  reg        [376:0]  stage1_inputData_0_delay_32_X;
  reg        [376:0]  stage1_inputData_0_delay_32_Y;
  reg        [376:0]  stage1_inputData_0_delay_32_Z;
  reg        [376:0]  stage1_inputData_0_delay_32_T;
  reg        [376:0]  stage1_inputData_0_delay_33_X;
  reg        [376:0]  stage1_inputData_0_delay_33_Y;
  reg        [376:0]  stage1_inputData_0_delay_33_Z;
  reg        [376:0]  stage1_inputData_0_delay_33_T;
  reg        [376:0]  stage1_inputData_0_delay_34_X;
  reg        [376:0]  stage1_inputData_0_delay_34_Y;
  reg        [376:0]  stage1_inputData_0_delay_34_Z;
  reg        [376:0]  stage1_inputData_0_delay_34_T;
  reg        [376:0]  stage1_inputData_0_delay_35_X;
  reg        [376:0]  stage1_inputData_0_delay_35_Y;
  reg        [376:0]  stage1_inputData_0_delay_35_Z;
  reg        [376:0]  stage1_inputData_0_delay_35_T;
  reg        [376:0]  pAddPort_0_s_delay_1_X;
  reg        [376:0]  pAddPort_0_s_delay_1_Y;
  reg        [376:0]  pAddPort_0_s_delay_1_Z;
  reg        [376:0]  pAddPort_0_s_delay_1_T;
  reg        [376:0]  pAddPort_0_s_delay_2_X;
  reg        [376:0]  pAddPort_0_s_delay_2_Y;
  reg        [376:0]  pAddPort_0_s_delay_2_Z;
  reg        [376:0]  pAddPort_0_s_delay_2_T;
  reg        [376:0]  pAddPort_0_s_delay_3_X;
  reg        [376:0]  pAddPort_0_s_delay_3_Y;
  reg        [376:0]  pAddPort_0_s_delay_3_Z;
  reg        [376:0]  pAddPort_0_s_delay_3_T;
  reg        [376:0]  pAddPort_0_s_delay_4_X;
  reg        [376:0]  pAddPort_0_s_delay_4_Y;
  reg        [376:0]  pAddPort_0_s_delay_4_Z;
  reg        [376:0]  pAddPort_0_s_delay_4_T;
  reg        [376:0]  pAddPort_0_s_delay_5_X;
  reg        [376:0]  pAddPort_0_s_delay_5_Y;
  reg        [376:0]  pAddPort_0_s_delay_5_Z;
  reg        [376:0]  pAddPort_0_s_delay_5_T;
  reg        [376:0]  pAddPort_0_s_delay_6_X;
  reg        [376:0]  pAddPort_0_s_delay_6_Y;
  reg        [376:0]  pAddPort_0_s_delay_6_Z;
  reg        [376:0]  pAddPort_0_s_delay_6_T;
  reg        [376:0]  pAddPort_0_s_delay_7_X;
  reg        [376:0]  pAddPort_0_s_delay_7_Y;
  reg        [376:0]  pAddPort_0_s_delay_7_Z;
  reg        [376:0]  pAddPort_0_s_delay_7_T;
  reg        [376:0]  pAddPort_0_s_delay_8_X;
  reg        [376:0]  pAddPort_0_s_delay_8_Y;
  reg        [376:0]  pAddPort_0_s_delay_8_Z;
  reg        [376:0]  pAddPort_0_s_delay_8_T;
  reg        [376:0]  pAddPort_0_s_delay_9_X;
  reg        [376:0]  pAddPort_0_s_delay_9_Y;
  reg        [376:0]  pAddPort_0_s_delay_9_Z;
  reg        [376:0]  pAddPort_0_s_delay_9_T;
  reg        [376:0]  pAddPort_0_s_delay_10_X;
  reg        [376:0]  pAddPort_0_s_delay_10_Y;
  reg        [376:0]  pAddPort_0_s_delay_10_Z;
  reg        [376:0]  pAddPort_0_s_delay_10_T;
  reg        [376:0]  pAddPort_0_s_delay_11_X;
  reg        [376:0]  pAddPort_0_s_delay_11_Y;
  reg        [376:0]  pAddPort_0_s_delay_11_Z;
  reg        [376:0]  pAddPort_0_s_delay_11_T;
  reg        [376:0]  pAddPort_0_s_delay_12_X;
  reg        [376:0]  pAddPort_0_s_delay_12_Y;
  reg        [376:0]  pAddPort_0_s_delay_12_Z;
  reg        [376:0]  pAddPort_0_s_delay_12_T;
  reg        [376:0]  pAddPort_0_s_delay_13_X;
  reg        [376:0]  pAddPort_0_s_delay_13_Y;
  reg        [376:0]  pAddPort_0_s_delay_13_Z;
  reg        [376:0]  pAddPort_0_s_delay_13_T;
  reg        [376:0]  pAddPort_0_s_delay_14_X;
  reg        [376:0]  pAddPort_0_s_delay_14_Y;
  reg        [376:0]  pAddPort_0_s_delay_14_Z;
  reg        [376:0]  pAddPort_0_s_delay_14_T;
  reg        [376:0]  pAddPort_0_s_delay_15_X;
  reg        [376:0]  pAddPort_0_s_delay_15_Y;
  reg        [376:0]  pAddPort_0_s_delay_15_Z;
  reg        [376:0]  pAddPort_0_s_delay_15_T;
  reg        [376:0]  pAddPort_0_s_delay_16_X;
  reg        [376:0]  pAddPort_0_s_delay_16_Y;
  reg        [376:0]  pAddPort_0_s_delay_16_Z;
  reg        [376:0]  pAddPort_0_s_delay_16_T;
  reg        [376:0]  pAddPort_0_s_delay_17_X;
  reg        [376:0]  pAddPort_0_s_delay_17_Y;
  reg        [376:0]  pAddPort_0_s_delay_17_Z;
  reg        [376:0]  pAddPort_0_s_delay_17_T;
  reg        [376:0]  pAddPort_0_s_delay_18_X;
  reg        [376:0]  pAddPort_0_s_delay_18_Y;
  reg        [376:0]  pAddPort_0_s_delay_18_Z;
  reg        [376:0]  pAddPort_0_s_delay_18_T;
  reg        [376:0]  pAddPort_0_s_delay_19_X;
  reg        [376:0]  pAddPort_0_s_delay_19_Y;
  reg        [376:0]  pAddPort_0_s_delay_19_Z;
  reg        [376:0]  pAddPort_0_s_delay_19_T;
  reg        [376:0]  pAddPort_0_s_delay_20_X;
  reg        [376:0]  pAddPort_0_s_delay_20_Y;
  reg        [376:0]  pAddPort_0_s_delay_20_Z;
  reg        [376:0]  pAddPort_0_s_delay_20_T;
  reg        [376:0]  pAddPort_0_s_delay_21_X;
  reg        [376:0]  pAddPort_0_s_delay_21_Y;
  reg        [376:0]  pAddPort_0_s_delay_21_Z;
  reg        [376:0]  pAddPort_0_s_delay_21_T;
  reg        [376:0]  pAddPort_0_s_delay_22_X;
  reg        [376:0]  pAddPort_0_s_delay_22_Y;
  reg        [376:0]  pAddPort_0_s_delay_22_Z;
  reg        [376:0]  pAddPort_0_s_delay_22_T;
  reg        [376:0]  pAddPort_0_s_delay_23_X;
  reg        [376:0]  pAddPort_0_s_delay_23_Y;
  reg        [376:0]  pAddPort_0_s_delay_23_Z;
  reg        [376:0]  pAddPort_0_s_delay_23_T;
  reg        [376:0]  pAddPort_0_s_delay_24_X;
  reg        [376:0]  pAddPort_0_s_delay_24_Y;
  reg        [376:0]  pAddPort_0_s_delay_24_Z;
  reg        [376:0]  pAddPort_0_s_delay_24_T;
  reg        [376:0]  pAddPort_0_s_delay_25_X;
  reg        [376:0]  pAddPort_0_s_delay_25_Y;
  reg        [376:0]  pAddPort_0_s_delay_25_Z;
  reg        [376:0]  pAddPort_0_s_delay_25_T;
  reg        [376:0]  pAddPort_0_s_delay_26_X;
  reg        [376:0]  pAddPort_0_s_delay_26_Y;
  reg        [376:0]  pAddPort_0_s_delay_26_Z;
  reg        [376:0]  pAddPort_0_s_delay_26_T;
  reg        [376:0]  pAddPort_0_s_delay_27_X;
  reg        [376:0]  pAddPort_0_s_delay_27_Y;
  reg        [376:0]  pAddPort_0_s_delay_27_Z;
  reg        [376:0]  pAddPort_0_s_delay_27_T;
  reg        [376:0]  pAddPort_0_s_delay_28_X;
  reg        [376:0]  pAddPort_0_s_delay_28_Y;
  reg        [376:0]  pAddPort_0_s_delay_28_Z;
  reg        [376:0]  pAddPort_0_s_delay_28_T;
  reg        [376:0]  pAddPort_0_s_delay_29_X;
  reg        [376:0]  pAddPort_0_s_delay_29_Y;
  reg        [376:0]  pAddPort_0_s_delay_29_Z;
  reg        [376:0]  pAddPort_0_s_delay_29_T;
  reg        [376:0]  pAddPort_0_s_delay_30_X;
  reg        [376:0]  pAddPort_0_s_delay_30_Y;
  reg        [376:0]  pAddPort_0_s_delay_30_Z;
  reg        [376:0]  pAddPort_0_s_delay_30_T;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_1;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_2;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_3;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_4;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_5;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_6;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_7;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_8;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_9;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_10;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_11;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_12;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_13;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_14;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_15;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_16;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_17;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_18;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_19;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_20;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_21;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_22;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_23;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_24;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_25;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_26;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_27;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_28;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_29;
  reg        [15:0]   shiftRegs_addressOutFull_0_delay_30;
  reg                 _zz_io_dataIn_1_valid;
  reg                 _zz_io_dataIn_1_valid_1;
  reg                 _zz_io_dataIn_1_valid_2;
  reg                 _zz_io_dataIn_1_valid_3;
  reg                 _zz_io_dataIn_1_valid_4;
  reg                 _zz_io_dataIn_1_valid_5;
  reg                 _zz_io_dataIn_1_valid_6;
  reg                 _zz_io_dataIn_1_valid_7;
  reg                 _zz_io_dataIn_1_valid_8;
  reg                 _zz_io_dataIn_1_valid_9;
  reg                 _zz_io_dataIn_1_valid_10;
  reg                 _zz_io_dataIn_1_valid_11;
  reg                 _zz_io_dataIn_1_valid_12;
  reg                 _zz_io_dataIn_1_valid_13;
  reg                 _zz_io_dataIn_1_valid_14;
  reg                 _zz_io_dataIn_1_valid_15;
  reg                 _zz_io_dataIn_1_valid_16;
  reg                 _zz_io_dataIn_1_valid_17;
  reg                 _zz_io_dataIn_1_valid_18;
  reg                 _zz_io_dataIn_1_valid_19;
  reg                 _zz_io_dataIn_1_valid_20;
  reg                 _zz_io_dataIn_1_valid_21;
  reg                 _zz_io_dataIn_1_valid_22;
  reg                 _zz_io_dataIn_1_valid_23;
  reg                 _zz_io_dataIn_1_valid_24;
  reg                 _zz_io_dataIn_1_valid_25;
  reg                 _zz_io_dataIn_1_valid_26;
  reg                 _zz_io_dataIn_1_valid_27;
  reg                 _zz_io_dataIn_1_valid_28;
  reg                 _zz_io_dataIn_1_valid_29;
  reg                 _zz_io_dataIn_1_valid_30;
  reg                 _zz_io_dataIn_1_valid_31;
  reg                 _zz_io_dataIn_1_valid_32;
  reg                 _zz_io_dataIn_1_valid_33;
  reg                 _zz_io_dataIn_1_valid_34;
  reg        [376:0]  stage1_inputData_0_delay_1_X_2;
  reg        [376:0]  stage1_inputData_0_delay_1_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_1_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_1_T_2;
  reg        [376:0]  stage1_inputData_0_delay_2_X_2;
  reg        [376:0]  stage1_inputData_0_delay_2_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_2_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_2_T_2;
  reg        [376:0]  stage1_inputData_0_delay_3_X_2;
  reg        [376:0]  stage1_inputData_0_delay_3_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_3_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_3_T_2;
  reg        [376:0]  stage1_inputData_0_delay_4_X_2;
  reg        [376:0]  stage1_inputData_0_delay_4_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_4_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_4_T_2;
  reg        [376:0]  stage1_inputData_0_delay_5_X_2;
  reg        [376:0]  stage1_inputData_0_delay_5_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_5_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_5_T_2;
  reg        [376:0]  stage1_inputData_0_delay_6_X_1;
  reg        [376:0]  stage1_inputData_0_delay_6_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_6_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_6_T_1;
  reg        [376:0]  stage1_inputData_0_delay_7_X_1;
  reg        [376:0]  stage1_inputData_0_delay_7_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_7_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_7_T_1;
  reg        [376:0]  stage1_inputData_0_delay_8_X_1;
  reg        [376:0]  stage1_inputData_0_delay_8_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_8_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_8_T_1;
  reg        [376:0]  stage1_inputData_0_delay_9_X_1;
  reg        [376:0]  stage1_inputData_0_delay_9_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_9_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_9_T_1;
  reg        [376:0]  stage1_inputData_0_delay_10_X_1;
  reg        [376:0]  stage1_inputData_0_delay_10_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_10_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_10_T_1;
  reg        [376:0]  stage1_inputData_0_delay_11_X_1;
  reg        [376:0]  stage1_inputData_0_delay_11_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_11_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_11_T_1;
  reg        [376:0]  stage1_inputData_0_delay_12_X_1;
  reg        [376:0]  stage1_inputData_0_delay_12_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_12_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_12_T_1;
  reg        [376:0]  stage1_inputData_0_delay_13_X_1;
  reg        [376:0]  stage1_inputData_0_delay_13_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_13_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_13_T_1;
  reg        [376:0]  stage1_inputData_0_delay_14_X_1;
  reg        [376:0]  stage1_inputData_0_delay_14_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_14_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_14_T_1;
  reg        [376:0]  stage1_inputData_0_delay_15_X_1;
  reg        [376:0]  stage1_inputData_0_delay_15_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_15_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_15_T_1;
  reg        [376:0]  stage1_inputData_0_delay_16_X_1;
  reg        [376:0]  stage1_inputData_0_delay_16_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_16_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_16_T_1;
  reg        [376:0]  stage1_inputData_0_delay_17_X_1;
  reg        [376:0]  stage1_inputData_0_delay_17_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_17_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_17_T_1;
  reg        [376:0]  stage1_inputData_0_delay_18_X_1;
  reg        [376:0]  stage1_inputData_0_delay_18_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_18_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_18_T_1;
  reg        [376:0]  stage1_inputData_0_delay_19_X_1;
  reg        [376:0]  stage1_inputData_0_delay_19_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_19_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_19_T_1;
  reg        [376:0]  stage1_inputData_0_delay_20_X_1;
  reg        [376:0]  stage1_inputData_0_delay_20_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_20_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_20_T_1;
  reg        [376:0]  stage1_inputData_0_delay_21_X_1;
  reg        [376:0]  stage1_inputData_0_delay_21_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_21_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_21_T_1;
  reg        [376:0]  stage1_inputData_0_delay_22_X_1;
  reg        [376:0]  stage1_inputData_0_delay_22_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_22_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_22_T_1;
  reg        [376:0]  stage1_inputData_0_delay_23_X_1;
  reg        [376:0]  stage1_inputData_0_delay_23_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_23_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_23_T_1;
  reg        [376:0]  stage1_inputData_0_delay_24_X_1;
  reg        [376:0]  stage1_inputData_0_delay_24_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_24_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_24_T_1;
  reg        [376:0]  stage1_inputData_0_delay_25_X_1;
  reg        [376:0]  stage1_inputData_0_delay_25_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_25_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_25_T_1;
  reg        [376:0]  stage1_inputData_0_delay_26_X_1;
  reg        [376:0]  stage1_inputData_0_delay_26_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_26_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_26_T_1;
  reg        [376:0]  stage1_inputData_0_delay_27_X_1;
  reg        [376:0]  stage1_inputData_0_delay_27_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_27_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_27_T_1;
  reg        [376:0]  stage1_inputData_0_delay_28_X_1;
  reg        [376:0]  stage1_inputData_0_delay_28_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_28_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_28_T_1;
  reg        [376:0]  stage1_inputData_0_delay_29_X_1;
  reg        [376:0]  stage1_inputData_0_delay_29_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_29_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_29_T_1;
  reg        [376:0]  stage1_inputData_0_delay_30_X_1;
  reg        [376:0]  stage1_inputData_0_delay_30_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_30_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_30_T_1;
  reg        [376:0]  stage1_inputData_0_delay_31_X_1;
  reg        [376:0]  stage1_inputData_0_delay_31_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_31_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_31_T_1;
  reg        [376:0]  stage1_inputData_0_delay_32_X_1;
  reg        [376:0]  stage1_inputData_0_delay_32_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_32_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_32_T_1;
  reg        [376:0]  stage1_inputData_0_delay_33_X_1;
  reg        [376:0]  stage1_inputData_0_delay_33_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_33_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_33_T_1;
  reg        [376:0]  stage1_inputData_0_delay_34_X_1;
  reg        [376:0]  stage1_inputData_0_delay_34_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_34_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_34_T_1;
  reg        [376:0]  stage1_inputData_0_delay_35_X_1;
  reg        [376:0]  stage1_inputData_0_delay_35_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_35_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_35_T_1;
  reg        [15:0]   stage1_inputAddress_0_delay_1_1;
  reg        [15:0]   stage1_inputAddress_0_delay_2_1;
  reg        [15:0]   stage1_inputAddress_0_delay_3_1;
  reg        [15:0]   stage1_inputAddress_0_delay_4_1;
  reg        [15:0]   stage1_inputAddress_0_delay_5_1;
  reg        [15:0]   stage1_inputAddress_0_delay_6;
  reg        [15:0]   stage1_inputAddress_0_delay_7;
  reg        [15:0]   stage1_inputAddress_0_delay_8;
  reg        [15:0]   stage1_inputAddress_0_delay_9;
  reg        [15:0]   stage1_inputAddress_0_delay_10;
  reg        [15:0]   stage1_inputAddress_0_delay_11;
  reg        [15:0]   stage1_inputAddress_0_delay_12;
  reg        [15:0]   stage1_inputAddress_0_delay_13;
  reg        [15:0]   stage1_inputAddress_0_delay_14;
  reg        [15:0]   stage1_inputAddress_0_delay_15;
  reg        [15:0]   stage1_inputAddress_0_delay_16;
  reg        [15:0]   stage1_inputAddress_0_delay_17;
  reg        [15:0]   stage1_inputAddress_0_delay_18;
  reg        [15:0]   stage1_inputAddress_0_delay_19;
  reg        [15:0]   stage1_inputAddress_0_delay_20;
  reg        [15:0]   stage1_inputAddress_0_delay_21;
  reg        [15:0]   stage1_inputAddress_0_delay_22;
  reg        [15:0]   stage1_inputAddress_0_delay_23;
  reg        [15:0]   stage1_inputAddress_0_delay_24;
  reg        [15:0]   stage1_inputAddress_0_delay_25;
  reg        [15:0]   stage1_inputAddress_0_delay_26;
  reg        [15:0]   stage1_inputAddress_0_delay_27;
  reg        [15:0]   stage1_inputAddress_0_delay_28;
  reg        [15:0]   stage1_inputAddress_0_delay_29;
  reg        [15:0]   stage1_inputAddress_0_delay_30;
  reg        [15:0]   stage1_inputAddress_0_delay_31;
  reg        [15:0]   stage1_inputAddress_0_delay_32;
  reg        [15:0]   stage1_inputAddress_0_delay_33;
  reg        [15:0]   stage1_inputAddress_0_delay_34;
  reg        [15:0]   stage1_inputAddress_0_delay_35;
  reg                 stage1_inputValid_1_delay_1;
  reg                 stage1_inputValid_1_delay_2;
  reg                 stage1_inputValid_1_delay_3;
  reg                 stage1_inputValid_1_delay_4;
  reg                 stage1_inputValid_1_delay_5;
  reg        [15:0]   stage1_inputAddress_1_delay_1;
  reg        [15:0]   stage1_inputAddress_1_delay_2;
  reg        [15:0]   stage1_inputAddress_1_delay_3;
  reg        [15:0]   stage1_inputAddress_1_delay_4;
  reg        [15:0]   stage1_inputAddress_1_delay_5;
  reg        [376:0]  stage1_inputData_1_delay_1_X;
  reg        [376:0]  stage1_inputData_1_delay_1_Y;
  reg        [376:0]  stage1_inputData_1_delay_1_Z;
  reg        [376:0]  stage1_inputData_1_delay_1_T;
  reg        [376:0]  stage1_inputData_1_delay_2_X;
  reg        [376:0]  stage1_inputData_1_delay_2_Y;
  reg        [376:0]  stage1_inputData_1_delay_2_Z;
  reg        [376:0]  stage1_inputData_1_delay_2_T;
  reg        [376:0]  stage1_inputData_1_delay_3_X;
  reg        [376:0]  stage1_inputData_1_delay_3_Y;
  reg        [376:0]  stage1_inputData_1_delay_3_Z;
  reg        [376:0]  stage1_inputData_1_delay_3_T;
  reg        [376:0]  stage1_inputData_1_delay_4_X;
  reg        [376:0]  stage1_inputData_1_delay_4_Y;
  reg        [376:0]  stage1_inputData_1_delay_4_Z;
  reg        [376:0]  stage1_inputData_1_delay_4_T;
  reg        [376:0]  stage1_inputData_1_delay_5_X;
  reg        [376:0]  stage1_inputData_1_delay_5_Y;
  reg        [376:0]  stage1_inputData_1_delay_5_Z;
  reg        [376:0]  stage1_inputData_1_delay_5_T;
  reg                 _zz_io_dataIn_0_valid_35;
  reg                 _zz_io_dataIn_0_valid_36;
  reg                 _zz_io_dataIn_0_valid_37;
  reg                 _zz_io_dataIn_0_valid_38;
  reg                 _zz_io_dataIn_0_valid_39;
  reg                 _zz_io_dataIn_0_valid_40;
  reg                 _zz_io_dataIn_0_valid_41;
  reg                 _zz_io_dataIn_0_valid_42;
  reg                 _zz_io_dataIn_0_valid_43;
  reg                 _zz_io_dataIn_0_valid_44;
  reg                 _zz_io_dataIn_0_valid_45;
  reg                 _zz_io_dataIn_0_valid_46;
  reg                 _zz_io_dataIn_0_valid_47;
  reg                 _zz_io_dataIn_0_valid_48;
  reg                 _zz_io_dataIn_0_valid_49;
  reg                 _zz_io_dataIn_0_valid_50;
  reg                 _zz_io_dataIn_0_valid_51;
  reg                 _zz_io_dataIn_0_valid_52;
  reg                 _zz_io_dataIn_0_valid_53;
  reg                 _zz_io_dataIn_0_valid_54;
  reg                 _zz_io_dataIn_0_valid_55;
  reg                 _zz_io_dataIn_0_valid_56;
  reg                 _zz_io_dataIn_0_valid_57;
  reg                 _zz_io_dataIn_0_valid_58;
  reg                 _zz_io_dataIn_0_valid_59;
  reg                 _zz_io_dataIn_0_valid_60;
  reg                 _zz_io_dataIn_0_valid_61;
  reg                 _zz_io_dataIn_0_valid_62;
  reg                 _zz_io_dataIn_0_valid_63;
  reg                 _zz_io_dataIn_0_valid_64;
  reg                 _zz_io_dataIn_0_valid_65;
  reg                 _zz_io_dataIn_0_valid_66;
  reg                 _zz_io_dataIn_0_valid_67;
  reg                 _zz_io_dataIn_0_valid_68;
  reg                 _zz_io_dataIn_0_valid_69;
  reg                 _zz_io_dataIn_0_payload_a_X_35;
  reg                 _zz_io_dataIn_0_payload_a_X_36;
  reg                 _zz_io_dataIn_0_payload_a_X_37;
  reg                 _zz_io_dataIn_0_payload_a_X_38;
  reg                 _zz_io_dataIn_0_payload_a_X_39;
  reg                 _zz_io_dataIn_0_payload_a_X_40;
  reg                 _zz_io_dataIn_0_payload_a_X_41;
  reg                 _zz_io_dataIn_0_payload_a_X_42;
  reg                 _zz_io_dataIn_0_payload_a_X_43;
  reg                 _zz_io_dataIn_0_payload_a_X_44;
  reg                 _zz_io_dataIn_0_payload_a_X_45;
  reg                 _zz_io_dataIn_0_payload_a_X_46;
  reg                 _zz_io_dataIn_0_payload_a_X_47;
  reg                 _zz_io_dataIn_0_payload_a_X_48;
  reg                 _zz_io_dataIn_0_payload_a_X_49;
  reg                 _zz_io_dataIn_0_payload_a_X_50;
  reg                 _zz_io_dataIn_0_payload_a_X_51;
  reg                 _zz_io_dataIn_0_payload_a_X_52;
  reg                 _zz_io_dataIn_0_payload_a_X_53;
  reg                 _zz_io_dataIn_0_payload_a_X_54;
  reg                 _zz_io_dataIn_0_payload_a_X_55;
  reg                 _zz_io_dataIn_0_payload_a_X_56;
  reg                 _zz_io_dataIn_0_payload_a_X_57;
  reg                 _zz_io_dataIn_0_payload_a_X_58;
  reg                 _zz_io_dataIn_0_payload_a_X_59;
  reg                 _zz_io_dataIn_0_payload_a_X_60;
  reg                 _zz_io_dataIn_0_payload_a_X_61;
  reg                 _zz_io_dataIn_0_payload_a_X_62;
  reg                 _zz_io_dataIn_0_payload_a_X_63;
  reg                 _zz_io_dataIn_0_payload_a_X_64;
  reg                 _zz_io_dataIn_0_payload_a_X_65;
  reg                 _zz_io_dataIn_0_payload_a_X_66;
  reg                 _zz_io_dataIn_0_payload_a_X_67;
  reg                 _zz_io_dataIn_0_payload_a_X_68;
  reg                 _zz_io_dataIn_0_payload_a_X_69;
  reg        [376:0]  stage1_inputData_1_delay_1_X_1;
  reg        [376:0]  stage1_inputData_1_delay_1_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_1_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_1_T_1;
  reg        [376:0]  stage1_inputData_1_delay_2_X_1;
  reg        [376:0]  stage1_inputData_1_delay_2_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_2_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_2_T_1;
  reg        [376:0]  stage1_inputData_1_delay_3_X_1;
  reg        [376:0]  stage1_inputData_1_delay_3_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_3_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_3_T_1;
  reg        [376:0]  stage1_inputData_1_delay_4_X_1;
  reg        [376:0]  stage1_inputData_1_delay_4_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_4_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_4_T_1;
  reg        [376:0]  stage1_inputData_1_delay_5_X_1;
  reg        [376:0]  stage1_inputData_1_delay_5_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_5_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_5_T_1;
  reg        [376:0]  stage1_inputData_1_delay_6_X;
  reg        [376:0]  stage1_inputData_1_delay_6_Y;
  reg        [376:0]  stage1_inputData_1_delay_6_Z;
  reg        [376:0]  stage1_inputData_1_delay_6_T;
  reg        [376:0]  stage1_inputData_1_delay_7_X;
  reg        [376:0]  stage1_inputData_1_delay_7_Y;
  reg        [376:0]  stage1_inputData_1_delay_7_Z;
  reg        [376:0]  stage1_inputData_1_delay_7_T;
  reg        [376:0]  stage1_inputData_1_delay_8_X;
  reg        [376:0]  stage1_inputData_1_delay_8_Y;
  reg        [376:0]  stage1_inputData_1_delay_8_Z;
  reg        [376:0]  stage1_inputData_1_delay_8_T;
  reg        [376:0]  stage1_inputData_1_delay_9_X;
  reg        [376:0]  stage1_inputData_1_delay_9_Y;
  reg        [376:0]  stage1_inputData_1_delay_9_Z;
  reg        [376:0]  stage1_inputData_1_delay_9_T;
  reg        [376:0]  stage1_inputData_1_delay_10_X;
  reg        [376:0]  stage1_inputData_1_delay_10_Y;
  reg        [376:0]  stage1_inputData_1_delay_10_Z;
  reg        [376:0]  stage1_inputData_1_delay_10_T;
  reg        [376:0]  stage1_inputData_1_delay_11_X;
  reg        [376:0]  stage1_inputData_1_delay_11_Y;
  reg        [376:0]  stage1_inputData_1_delay_11_Z;
  reg        [376:0]  stage1_inputData_1_delay_11_T;
  reg        [376:0]  stage1_inputData_1_delay_12_X;
  reg        [376:0]  stage1_inputData_1_delay_12_Y;
  reg        [376:0]  stage1_inputData_1_delay_12_Z;
  reg        [376:0]  stage1_inputData_1_delay_12_T;
  reg        [376:0]  stage1_inputData_1_delay_13_X;
  reg        [376:0]  stage1_inputData_1_delay_13_Y;
  reg        [376:0]  stage1_inputData_1_delay_13_Z;
  reg        [376:0]  stage1_inputData_1_delay_13_T;
  reg        [376:0]  stage1_inputData_1_delay_14_X;
  reg        [376:0]  stage1_inputData_1_delay_14_Y;
  reg        [376:0]  stage1_inputData_1_delay_14_Z;
  reg        [376:0]  stage1_inputData_1_delay_14_T;
  reg        [376:0]  stage1_inputData_1_delay_15_X;
  reg        [376:0]  stage1_inputData_1_delay_15_Y;
  reg        [376:0]  stage1_inputData_1_delay_15_Z;
  reg        [376:0]  stage1_inputData_1_delay_15_T;
  reg        [376:0]  stage1_inputData_1_delay_16_X;
  reg        [376:0]  stage1_inputData_1_delay_16_Y;
  reg        [376:0]  stage1_inputData_1_delay_16_Z;
  reg        [376:0]  stage1_inputData_1_delay_16_T;
  reg        [376:0]  stage1_inputData_1_delay_17_X;
  reg        [376:0]  stage1_inputData_1_delay_17_Y;
  reg        [376:0]  stage1_inputData_1_delay_17_Z;
  reg        [376:0]  stage1_inputData_1_delay_17_T;
  reg        [376:0]  stage1_inputData_1_delay_18_X;
  reg        [376:0]  stage1_inputData_1_delay_18_Y;
  reg        [376:0]  stage1_inputData_1_delay_18_Z;
  reg        [376:0]  stage1_inputData_1_delay_18_T;
  reg        [376:0]  stage1_inputData_1_delay_19_X;
  reg        [376:0]  stage1_inputData_1_delay_19_Y;
  reg        [376:0]  stage1_inputData_1_delay_19_Z;
  reg        [376:0]  stage1_inputData_1_delay_19_T;
  reg        [376:0]  stage1_inputData_1_delay_20_X;
  reg        [376:0]  stage1_inputData_1_delay_20_Y;
  reg        [376:0]  stage1_inputData_1_delay_20_Z;
  reg        [376:0]  stage1_inputData_1_delay_20_T;
  reg        [376:0]  stage1_inputData_1_delay_21_X;
  reg        [376:0]  stage1_inputData_1_delay_21_Y;
  reg        [376:0]  stage1_inputData_1_delay_21_Z;
  reg        [376:0]  stage1_inputData_1_delay_21_T;
  reg        [376:0]  stage1_inputData_1_delay_22_X;
  reg        [376:0]  stage1_inputData_1_delay_22_Y;
  reg        [376:0]  stage1_inputData_1_delay_22_Z;
  reg        [376:0]  stage1_inputData_1_delay_22_T;
  reg        [376:0]  stage1_inputData_1_delay_23_X;
  reg        [376:0]  stage1_inputData_1_delay_23_Y;
  reg        [376:0]  stage1_inputData_1_delay_23_Z;
  reg        [376:0]  stage1_inputData_1_delay_23_T;
  reg        [376:0]  stage1_inputData_1_delay_24_X;
  reg        [376:0]  stage1_inputData_1_delay_24_Y;
  reg        [376:0]  stage1_inputData_1_delay_24_Z;
  reg        [376:0]  stage1_inputData_1_delay_24_T;
  reg        [376:0]  stage1_inputData_1_delay_25_X;
  reg        [376:0]  stage1_inputData_1_delay_25_Y;
  reg        [376:0]  stage1_inputData_1_delay_25_Z;
  reg        [376:0]  stage1_inputData_1_delay_25_T;
  reg        [376:0]  stage1_inputData_1_delay_26_X;
  reg        [376:0]  stage1_inputData_1_delay_26_Y;
  reg        [376:0]  stage1_inputData_1_delay_26_Z;
  reg        [376:0]  stage1_inputData_1_delay_26_T;
  reg        [376:0]  stage1_inputData_1_delay_27_X;
  reg        [376:0]  stage1_inputData_1_delay_27_Y;
  reg        [376:0]  stage1_inputData_1_delay_27_Z;
  reg        [376:0]  stage1_inputData_1_delay_27_T;
  reg        [376:0]  stage1_inputData_1_delay_28_X;
  reg        [376:0]  stage1_inputData_1_delay_28_Y;
  reg        [376:0]  stage1_inputData_1_delay_28_Z;
  reg        [376:0]  stage1_inputData_1_delay_28_T;
  reg        [376:0]  stage1_inputData_1_delay_29_X;
  reg        [376:0]  stage1_inputData_1_delay_29_Y;
  reg        [376:0]  stage1_inputData_1_delay_29_Z;
  reg        [376:0]  stage1_inputData_1_delay_29_T;
  reg        [376:0]  stage1_inputData_1_delay_30_X;
  reg        [376:0]  stage1_inputData_1_delay_30_Y;
  reg        [376:0]  stage1_inputData_1_delay_30_Z;
  reg        [376:0]  stage1_inputData_1_delay_30_T;
  reg        [376:0]  stage1_inputData_1_delay_31_X;
  reg        [376:0]  stage1_inputData_1_delay_31_Y;
  reg        [376:0]  stage1_inputData_1_delay_31_Z;
  reg        [376:0]  stage1_inputData_1_delay_31_T;
  reg        [376:0]  stage1_inputData_1_delay_32_X;
  reg        [376:0]  stage1_inputData_1_delay_32_Y;
  reg        [376:0]  stage1_inputData_1_delay_32_Z;
  reg        [376:0]  stage1_inputData_1_delay_32_T;
  reg        [376:0]  stage1_inputData_1_delay_33_X;
  reg        [376:0]  stage1_inputData_1_delay_33_Y;
  reg        [376:0]  stage1_inputData_1_delay_33_Z;
  reg        [376:0]  stage1_inputData_1_delay_33_T;
  reg        [376:0]  stage1_inputData_1_delay_34_X;
  reg        [376:0]  stage1_inputData_1_delay_34_Y;
  reg        [376:0]  stage1_inputData_1_delay_34_Z;
  reg        [376:0]  stage1_inputData_1_delay_34_T;
  reg        [376:0]  stage1_inputData_1_delay_35_X;
  reg        [376:0]  stage1_inputData_1_delay_35_Y;
  reg        [376:0]  stage1_inputData_1_delay_35_Z;
  reg        [376:0]  stage1_inputData_1_delay_35_T;
  reg        [376:0]  pAddPort_1_s_delay_1_X;
  reg        [376:0]  pAddPort_1_s_delay_1_Y;
  reg        [376:0]  pAddPort_1_s_delay_1_Z;
  reg        [376:0]  pAddPort_1_s_delay_1_T;
  reg        [376:0]  pAddPort_1_s_delay_2_X;
  reg        [376:0]  pAddPort_1_s_delay_2_Y;
  reg        [376:0]  pAddPort_1_s_delay_2_Z;
  reg        [376:0]  pAddPort_1_s_delay_2_T;
  reg        [376:0]  pAddPort_1_s_delay_3_X;
  reg        [376:0]  pAddPort_1_s_delay_3_Y;
  reg        [376:0]  pAddPort_1_s_delay_3_Z;
  reg        [376:0]  pAddPort_1_s_delay_3_T;
  reg        [376:0]  pAddPort_1_s_delay_4_X;
  reg        [376:0]  pAddPort_1_s_delay_4_Y;
  reg        [376:0]  pAddPort_1_s_delay_4_Z;
  reg        [376:0]  pAddPort_1_s_delay_4_T;
  reg        [376:0]  pAddPort_1_s_delay_5_X;
  reg        [376:0]  pAddPort_1_s_delay_5_Y;
  reg        [376:0]  pAddPort_1_s_delay_5_Z;
  reg        [376:0]  pAddPort_1_s_delay_5_T;
  reg        [376:0]  pAddPort_1_s_delay_6_X;
  reg        [376:0]  pAddPort_1_s_delay_6_Y;
  reg        [376:0]  pAddPort_1_s_delay_6_Z;
  reg        [376:0]  pAddPort_1_s_delay_6_T;
  reg        [376:0]  pAddPort_1_s_delay_7_X;
  reg        [376:0]  pAddPort_1_s_delay_7_Y;
  reg        [376:0]  pAddPort_1_s_delay_7_Z;
  reg        [376:0]  pAddPort_1_s_delay_7_T;
  reg        [376:0]  pAddPort_1_s_delay_8_X;
  reg        [376:0]  pAddPort_1_s_delay_8_Y;
  reg        [376:0]  pAddPort_1_s_delay_8_Z;
  reg        [376:0]  pAddPort_1_s_delay_8_T;
  reg        [376:0]  pAddPort_1_s_delay_9_X;
  reg        [376:0]  pAddPort_1_s_delay_9_Y;
  reg        [376:0]  pAddPort_1_s_delay_9_Z;
  reg        [376:0]  pAddPort_1_s_delay_9_T;
  reg        [376:0]  pAddPort_1_s_delay_10_X;
  reg        [376:0]  pAddPort_1_s_delay_10_Y;
  reg        [376:0]  pAddPort_1_s_delay_10_Z;
  reg        [376:0]  pAddPort_1_s_delay_10_T;
  reg        [376:0]  pAddPort_1_s_delay_11_X;
  reg        [376:0]  pAddPort_1_s_delay_11_Y;
  reg        [376:0]  pAddPort_1_s_delay_11_Z;
  reg        [376:0]  pAddPort_1_s_delay_11_T;
  reg        [376:0]  pAddPort_1_s_delay_12_X;
  reg        [376:0]  pAddPort_1_s_delay_12_Y;
  reg        [376:0]  pAddPort_1_s_delay_12_Z;
  reg        [376:0]  pAddPort_1_s_delay_12_T;
  reg        [376:0]  pAddPort_1_s_delay_13_X;
  reg        [376:0]  pAddPort_1_s_delay_13_Y;
  reg        [376:0]  pAddPort_1_s_delay_13_Z;
  reg        [376:0]  pAddPort_1_s_delay_13_T;
  reg        [376:0]  pAddPort_1_s_delay_14_X;
  reg        [376:0]  pAddPort_1_s_delay_14_Y;
  reg        [376:0]  pAddPort_1_s_delay_14_Z;
  reg        [376:0]  pAddPort_1_s_delay_14_T;
  reg        [376:0]  pAddPort_1_s_delay_15_X;
  reg        [376:0]  pAddPort_1_s_delay_15_Y;
  reg        [376:0]  pAddPort_1_s_delay_15_Z;
  reg        [376:0]  pAddPort_1_s_delay_15_T;
  reg        [376:0]  pAddPort_1_s_delay_16_X;
  reg        [376:0]  pAddPort_1_s_delay_16_Y;
  reg        [376:0]  pAddPort_1_s_delay_16_Z;
  reg        [376:0]  pAddPort_1_s_delay_16_T;
  reg        [376:0]  pAddPort_1_s_delay_17_X;
  reg        [376:0]  pAddPort_1_s_delay_17_Y;
  reg        [376:0]  pAddPort_1_s_delay_17_Z;
  reg        [376:0]  pAddPort_1_s_delay_17_T;
  reg        [376:0]  pAddPort_1_s_delay_18_X;
  reg        [376:0]  pAddPort_1_s_delay_18_Y;
  reg        [376:0]  pAddPort_1_s_delay_18_Z;
  reg        [376:0]  pAddPort_1_s_delay_18_T;
  reg        [376:0]  pAddPort_1_s_delay_19_X;
  reg        [376:0]  pAddPort_1_s_delay_19_Y;
  reg        [376:0]  pAddPort_1_s_delay_19_Z;
  reg        [376:0]  pAddPort_1_s_delay_19_T;
  reg        [376:0]  pAddPort_1_s_delay_20_X;
  reg        [376:0]  pAddPort_1_s_delay_20_Y;
  reg        [376:0]  pAddPort_1_s_delay_20_Z;
  reg        [376:0]  pAddPort_1_s_delay_20_T;
  reg        [376:0]  pAddPort_1_s_delay_21_X;
  reg        [376:0]  pAddPort_1_s_delay_21_Y;
  reg        [376:0]  pAddPort_1_s_delay_21_Z;
  reg        [376:0]  pAddPort_1_s_delay_21_T;
  reg        [376:0]  pAddPort_1_s_delay_22_X;
  reg        [376:0]  pAddPort_1_s_delay_22_Y;
  reg        [376:0]  pAddPort_1_s_delay_22_Z;
  reg        [376:0]  pAddPort_1_s_delay_22_T;
  reg        [376:0]  pAddPort_1_s_delay_23_X;
  reg        [376:0]  pAddPort_1_s_delay_23_Y;
  reg        [376:0]  pAddPort_1_s_delay_23_Z;
  reg        [376:0]  pAddPort_1_s_delay_23_T;
  reg        [376:0]  pAddPort_1_s_delay_24_X;
  reg        [376:0]  pAddPort_1_s_delay_24_Y;
  reg        [376:0]  pAddPort_1_s_delay_24_Z;
  reg        [376:0]  pAddPort_1_s_delay_24_T;
  reg        [376:0]  pAddPort_1_s_delay_25_X;
  reg        [376:0]  pAddPort_1_s_delay_25_Y;
  reg        [376:0]  pAddPort_1_s_delay_25_Z;
  reg        [376:0]  pAddPort_1_s_delay_25_T;
  reg        [376:0]  pAddPort_1_s_delay_26_X;
  reg        [376:0]  pAddPort_1_s_delay_26_Y;
  reg        [376:0]  pAddPort_1_s_delay_26_Z;
  reg        [376:0]  pAddPort_1_s_delay_26_T;
  reg        [376:0]  pAddPort_1_s_delay_27_X;
  reg        [376:0]  pAddPort_1_s_delay_27_Y;
  reg        [376:0]  pAddPort_1_s_delay_27_Z;
  reg        [376:0]  pAddPort_1_s_delay_27_T;
  reg        [376:0]  pAddPort_1_s_delay_28_X;
  reg        [376:0]  pAddPort_1_s_delay_28_Y;
  reg        [376:0]  pAddPort_1_s_delay_28_Z;
  reg        [376:0]  pAddPort_1_s_delay_28_T;
  reg        [376:0]  pAddPort_1_s_delay_29_X;
  reg        [376:0]  pAddPort_1_s_delay_29_Y;
  reg        [376:0]  pAddPort_1_s_delay_29_Z;
  reg        [376:0]  pAddPort_1_s_delay_29_T;
  reg        [376:0]  pAddPort_1_s_delay_30_X;
  reg        [376:0]  pAddPort_1_s_delay_30_Y;
  reg        [376:0]  pAddPort_1_s_delay_30_Z;
  reg        [376:0]  pAddPort_1_s_delay_30_T;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_1;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_2;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_3;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_4;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_5;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_6;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_7;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_8;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_9;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_10;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_11;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_12;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_13;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_14;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_15;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_16;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_17;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_18;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_19;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_20;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_21;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_22;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_23;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_24;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_25;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_26;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_27;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_28;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_29;
  reg        [15:0]   shiftRegs_addressOutFull_1_delay_30;
  reg                 _zz_io_dataIn_1_valid_35;
  reg                 _zz_io_dataIn_1_valid_36;
  reg                 _zz_io_dataIn_1_valid_37;
  reg                 _zz_io_dataIn_1_valid_38;
  reg                 _zz_io_dataIn_1_valid_39;
  reg                 _zz_io_dataIn_1_valid_40;
  reg                 _zz_io_dataIn_1_valid_41;
  reg                 _zz_io_dataIn_1_valid_42;
  reg                 _zz_io_dataIn_1_valid_43;
  reg                 _zz_io_dataIn_1_valid_44;
  reg                 _zz_io_dataIn_1_valid_45;
  reg                 _zz_io_dataIn_1_valid_46;
  reg                 _zz_io_dataIn_1_valid_47;
  reg                 _zz_io_dataIn_1_valid_48;
  reg                 _zz_io_dataIn_1_valid_49;
  reg                 _zz_io_dataIn_1_valid_50;
  reg                 _zz_io_dataIn_1_valid_51;
  reg                 _zz_io_dataIn_1_valid_52;
  reg                 _zz_io_dataIn_1_valid_53;
  reg                 _zz_io_dataIn_1_valid_54;
  reg                 _zz_io_dataIn_1_valid_55;
  reg                 _zz_io_dataIn_1_valid_56;
  reg                 _zz_io_dataIn_1_valid_57;
  reg                 _zz_io_dataIn_1_valid_58;
  reg                 _zz_io_dataIn_1_valid_59;
  reg                 _zz_io_dataIn_1_valid_60;
  reg                 _zz_io_dataIn_1_valid_61;
  reg                 _zz_io_dataIn_1_valid_62;
  reg                 _zz_io_dataIn_1_valid_63;
  reg                 _zz_io_dataIn_1_valid_64;
  reg                 _zz_io_dataIn_1_valid_65;
  reg                 _zz_io_dataIn_1_valid_66;
  reg                 _zz_io_dataIn_1_valid_67;
  reg                 _zz_io_dataIn_1_valid_68;
  reg                 _zz_io_dataIn_1_valid_69;
  reg        [376:0]  stage1_inputData_1_delay_1_X_2;
  reg        [376:0]  stage1_inputData_1_delay_1_Y_2;
  reg        [376:0]  stage1_inputData_1_delay_1_Z_2;
  reg        [376:0]  stage1_inputData_1_delay_1_T_2;
  reg        [376:0]  stage1_inputData_1_delay_2_X_2;
  reg        [376:0]  stage1_inputData_1_delay_2_Y_2;
  reg        [376:0]  stage1_inputData_1_delay_2_Z_2;
  reg        [376:0]  stage1_inputData_1_delay_2_T_2;
  reg        [376:0]  stage1_inputData_1_delay_3_X_2;
  reg        [376:0]  stage1_inputData_1_delay_3_Y_2;
  reg        [376:0]  stage1_inputData_1_delay_3_Z_2;
  reg        [376:0]  stage1_inputData_1_delay_3_T_2;
  reg        [376:0]  stage1_inputData_1_delay_4_X_2;
  reg        [376:0]  stage1_inputData_1_delay_4_Y_2;
  reg        [376:0]  stage1_inputData_1_delay_4_Z_2;
  reg        [376:0]  stage1_inputData_1_delay_4_T_2;
  reg        [376:0]  stage1_inputData_1_delay_5_X_2;
  reg        [376:0]  stage1_inputData_1_delay_5_Y_2;
  reg        [376:0]  stage1_inputData_1_delay_5_Z_2;
  reg        [376:0]  stage1_inputData_1_delay_5_T_2;
  reg        [376:0]  stage1_inputData_1_delay_6_X_1;
  reg        [376:0]  stage1_inputData_1_delay_6_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_6_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_6_T_1;
  reg        [376:0]  stage1_inputData_1_delay_7_X_1;
  reg        [376:0]  stage1_inputData_1_delay_7_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_7_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_7_T_1;
  reg        [376:0]  stage1_inputData_1_delay_8_X_1;
  reg        [376:0]  stage1_inputData_1_delay_8_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_8_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_8_T_1;
  reg        [376:0]  stage1_inputData_1_delay_9_X_1;
  reg        [376:0]  stage1_inputData_1_delay_9_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_9_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_9_T_1;
  reg        [376:0]  stage1_inputData_1_delay_10_X_1;
  reg        [376:0]  stage1_inputData_1_delay_10_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_10_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_10_T_1;
  reg        [376:0]  stage1_inputData_1_delay_11_X_1;
  reg        [376:0]  stage1_inputData_1_delay_11_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_11_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_11_T_1;
  reg        [376:0]  stage1_inputData_1_delay_12_X_1;
  reg        [376:0]  stage1_inputData_1_delay_12_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_12_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_12_T_1;
  reg        [376:0]  stage1_inputData_1_delay_13_X_1;
  reg        [376:0]  stage1_inputData_1_delay_13_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_13_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_13_T_1;
  reg        [376:0]  stage1_inputData_1_delay_14_X_1;
  reg        [376:0]  stage1_inputData_1_delay_14_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_14_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_14_T_1;
  reg        [376:0]  stage1_inputData_1_delay_15_X_1;
  reg        [376:0]  stage1_inputData_1_delay_15_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_15_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_15_T_1;
  reg        [376:0]  stage1_inputData_1_delay_16_X_1;
  reg        [376:0]  stage1_inputData_1_delay_16_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_16_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_16_T_1;
  reg        [376:0]  stage1_inputData_1_delay_17_X_1;
  reg        [376:0]  stage1_inputData_1_delay_17_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_17_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_17_T_1;
  reg        [376:0]  stage1_inputData_1_delay_18_X_1;
  reg        [376:0]  stage1_inputData_1_delay_18_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_18_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_18_T_1;
  reg        [376:0]  stage1_inputData_1_delay_19_X_1;
  reg        [376:0]  stage1_inputData_1_delay_19_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_19_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_19_T_1;
  reg        [376:0]  stage1_inputData_1_delay_20_X_1;
  reg        [376:0]  stage1_inputData_1_delay_20_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_20_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_20_T_1;
  reg        [376:0]  stage1_inputData_1_delay_21_X_1;
  reg        [376:0]  stage1_inputData_1_delay_21_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_21_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_21_T_1;
  reg        [376:0]  stage1_inputData_1_delay_22_X_1;
  reg        [376:0]  stage1_inputData_1_delay_22_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_22_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_22_T_1;
  reg        [376:0]  stage1_inputData_1_delay_23_X_1;
  reg        [376:0]  stage1_inputData_1_delay_23_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_23_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_23_T_1;
  reg        [376:0]  stage1_inputData_1_delay_24_X_1;
  reg        [376:0]  stage1_inputData_1_delay_24_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_24_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_24_T_1;
  reg        [376:0]  stage1_inputData_1_delay_25_X_1;
  reg        [376:0]  stage1_inputData_1_delay_25_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_25_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_25_T_1;
  reg        [376:0]  stage1_inputData_1_delay_26_X_1;
  reg        [376:0]  stage1_inputData_1_delay_26_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_26_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_26_T_1;
  reg        [376:0]  stage1_inputData_1_delay_27_X_1;
  reg        [376:0]  stage1_inputData_1_delay_27_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_27_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_27_T_1;
  reg        [376:0]  stage1_inputData_1_delay_28_X_1;
  reg        [376:0]  stage1_inputData_1_delay_28_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_28_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_28_T_1;
  reg        [376:0]  stage1_inputData_1_delay_29_X_1;
  reg        [376:0]  stage1_inputData_1_delay_29_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_29_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_29_T_1;
  reg        [376:0]  stage1_inputData_1_delay_30_X_1;
  reg        [376:0]  stage1_inputData_1_delay_30_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_30_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_30_T_1;
  reg        [376:0]  stage1_inputData_1_delay_31_X_1;
  reg        [376:0]  stage1_inputData_1_delay_31_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_31_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_31_T_1;
  reg        [376:0]  stage1_inputData_1_delay_32_X_1;
  reg        [376:0]  stage1_inputData_1_delay_32_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_32_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_32_T_1;
  reg        [376:0]  stage1_inputData_1_delay_33_X_1;
  reg        [376:0]  stage1_inputData_1_delay_33_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_33_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_33_T_1;
  reg        [376:0]  stage1_inputData_1_delay_34_X_1;
  reg        [376:0]  stage1_inputData_1_delay_34_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_34_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_34_T_1;
  reg        [376:0]  stage1_inputData_1_delay_35_X_1;
  reg        [376:0]  stage1_inputData_1_delay_35_Y_1;
  reg        [376:0]  stage1_inputData_1_delay_35_Z_1;
  reg        [376:0]  stage1_inputData_1_delay_35_T_1;
  reg        [15:0]   stage1_inputAddress_1_delay_1_1;
  reg        [15:0]   stage1_inputAddress_1_delay_2_1;
  reg        [15:0]   stage1_inputAddress_1_delay_3_1;
  reg        [15:0]   stage1_inputAddress_1_delay_4_1;
  reg        [15:0]   stage1_inputAddress_1_delay_5_1;
  reg        [15:0]   stage1_inputAddress_1_delay_6;
  reg        [15:0]   stage1_inputAddress_1_delay_7;
  reg        [15:0]   stage1_inputAddress_1_delay_8;
  reg        [15:0]   stage1_inputAddress_1_delay_9;
  reg        [15:0]   stage1_inputAddress_1_delay_10;
  reg        [15:0]   stage1_inputAddress_1_delay_11;
  reg        [15:0]   stage1_inputAddress_1_delay_12;
  reg        [15:0]   stage1_inputAddress_1_delay_13;
  reg        [15:0]   stage1_inputAddress_1_delay_14;
  reg        [15:0]   stage1_inputAddress_1_delay_15;
  reg        [15:0]   stage1_inputAddress_1_delay_16;
  reg        [15:0]   stage1_inputAddress_1_delay_17;
  reg        [15:0]   stage1_inputAddress_1_delay_18;
  reg        [15:0]   stage1_inputAddress_1_delay_19;
  reg        [15:0]   stage1_inputAddress_1_delay_20;
  reg        [15:0]   stage1_inputAddress_1_delay_21;
  reg        [15:0]   stage1_inputAddress_1_delay_22;
  reg        [15:0]   stage1_inputAddress_1_delay_23;
  reg        [15:0]   stage1_inputAddress_1_delay_24;
  reg        [15:0]   stage1_inputAddress_1_delay_25;
  reg        [15:0]   stage1_inputAddress_1_delay_26;
  reg        [15:0]   stage1_inputAddress_1_delay_27;
  reg        [15:0]   stage1_inputAddress_1_delay_28;
  reg        [15:0]   stage1_inputAddress_1_delay_29;
  reg        [15:0]   stage1_inputAddress_1_delay_30;
  reg        [15:0]   stage1_inputAddress_1_delay_31;
  reg        [15:0]   stage1_inputAddress_1_delay_32;
  reg        [15:0]   stage1_inputAddress_1_delay_33;
  reg        [15:0]   stage1_inputAddress_1_delay_34;
  reg        [15:0]   stage1_inputAddress_1_delay_35;
  wire                when_Pippenger_l153;
  wire                when_Pippenger_l168;
  reg                 _zz_io_state_1;
  reg                 _zz_io_state_1_1;
  reg                 _zz_io_state_1_2;
  reg                 _zz_io_state_1_3;
  reg                 _zz_io_state_1_4;
  reg                 _zz_io_state_1_5;
  reg                 _zz_io_state_1_6;
  reg                 _zz_io_state_1_7;
  reg                 _zz_io_state_1_8;
  reg                 _zz_io_state_1_9;
  reg                 _zz_io_state_1_10;
  reg                 _zz_io_state_1_11;
  reg                 _zz_io_state_1_12;
  reg                 _zz_io_state_1_13;
  reg                 _zz_io_state_1_14;
  reg                 _zz_io_state_1_15;
  reg                 _zz_io_state_1_16;
  reg                 _zz_io_state_1_17;
  reg                 _zz_io_state_1_18;
  reg                 _zz_io_state_1_19;
  reg                 _zz_io_state_1_20;
  reg                 _zz_io_state_1_21;
  reg                 _zz_io_state_1_22;
  reg                 _zz_io_state_1_23;
  reg                 _zz_io_state_1_24;
  reg                 _zz_io_state_1_25;
  reg                 _zz_io_state_1_26;
  reg                 _zz_io_state_1_27;
  reg                 _zz_io_state_1_28;
  reg                 _zz_io_state_1_29;
  reg                 _zz_io_state_1_30;
  reg                 _zz_io_state_1_31;
  reg                 _zz_io_state_1_32;
  reg                 _zz_io_state_1_33;
  reg                 _zz_io_state_1_34;
  reg                 _zz_io_state_1_35;
  reg                 _zz_io_state_1_36;
  reg                 _zz_io_state_1_37;
  reg                 _zz_io_state_1_38;
  reg                 _zz_io_dataIn_1_valid_70;
  reg                 _zz_io_dataIn_1_valid_71;
  reg                 _zz_io_dataIn_1_valid_72;
  reg                 _zz_io_dataIn_1_valid_73;
  reg                 _zz_io_dataIn_1_valid_74;
  reg                 _zz_io_dataIn_1_valid_75;
  reg                 _zz_io_dataIn_1_valid_76;
  reg                 _zz_io_dataIn_1_valid_77;
  reg                 _zz_io_dataIn_1_valid_78;
  reg                 _zz_io_dataIn_1_valid_79;
  reg                 _zz_io_dataIn_1_valid_80;
  reg                 _zz_io_dataIn_1_valid_81;
  reg                 _zz_io_dataIn_1_valid_82;
  reg                 _zz_io_dataIn_1_valid_83;
  reg                 _zz_io_dataIn_1_valid_84;
  reg                 _zz_io_dataIn_1_valid_85;
  reg                 _zz_io_dataIn_1_valid_86;
  reg                 _zz_io_dataIn_1_valid_87;
  reg                 _zz_io_dataIn_1_valid_88;
  reg                 _zz_io_dataIn_1_valid_89;
  reg                 _zz_io_dataIn_1_valid_90;
  reg                 _zz_io_dataIn_1_valid_91;
  reg                 _zz_io_dataIn_1_valid_92;
  reg                 _zz_io_dataIn_1_valid_93;
  reg                 _zz_io_dataIn_1_valid_94;
  reg                 _zz_io_dataIn_1_valid_95;
  reg                 _zz_io_dataIn_1_valid_96;
  reg                 _zz_io_dataIn_1_valid_97;
  reg                 _zz_io_dataIn_1_valid_98;
  reg                 _zz_io_dataIn_1_valid_99;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_X;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_Y;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_Z;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_T;
  reg        [15:0]   _zz_io_dataIn_1_payload_address;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_1;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_2;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_3;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_4;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_5;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_6;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_7;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_8;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_9;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_10;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_11;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_12;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_13;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_14;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_15;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_16;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_17;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_18;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_19;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_20;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_21;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_22;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_23;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_24;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_25;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_26;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_27;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_28;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_29;
  reg                 _zz_io_state_1_39;
  reg                 _zz_io_state_1_40;
  reg                 _zz_io_state_1_41;
  reg                 _zz_io_state_1_42;
  reg                 _zz_io_state_1_43;
  reg                 _zz_io_state_1_44;
  reg                 _zz_io_state_1_45;
  reg                 _zz_io_state_1_46;
  reg                 _zz_io_state_1_47;
  reg                 _zz_io_state_1_48;
  reg                 _zz_io_state_1_49;
  reg                 _zz_io_state_1_50;
  reg                 _zz_io_state_1_51;
  reg                 _zz_io_state_1_52;
  reg                 _zz_io_state_1_53;
  reg                 _zz_io_state_1_54;
  reg                 _zz_io_state_1_55;
  reg                 _zz_io_state_1_56;
  reg                 _zz_io_state_1_57;
  reg                 _zz_io_state_1_58;
  reg                 _zz_io_state_1_59;
  reg                 _zz_io_state_1_60;
  reg                 _zz_io_state_1_61;
  reg                 _zz_io_state_1_62;
  reg                 _zz_io_state_1_63;
  reg                 _zz_io_state_1_64;
  reg                 _zz_io_state_1_65;
  reg                 _zz_io_state_1_66;
  reg                 _zz_io_state_1_67;
  reg                 _zz_io_state_1_68;
  reg                 _zz_io_state_1_69;
  reg                 _zz_io_state_1_70;
  reg                 _zz_io_state_1_71;
  reg                 _zz_io_state_1_72;
  reg                 _zz_io_state_1_73;
  reg                 _zz_io_state_1_74;
  reg                 _zz_io_state_1_75;
  reg                 _zz_io_state_1_76;
  reg                 _zz_io_state_1_77;
  reg                 _zz_io_dataIn_1_valid_100;
  reg                 _zz_io_dataIn_1_valid_101;
  reg                 _zz_io_dataIn_1_valid_102;
  reg                 _zz_io_dataIn_1_valid_103;
  reg                 _zz_io_dataIn_1_valid_104;
  reg                 _zz_io_dataIn_1_valid_105;
  reg                 _zz_io_dataIn_1_valid_106;
  reg                 _zz_io_dataIn_1_valid_107;
  reg                 _zz_io_dataIn_1_valid_108;
  reg                 _zz_io_dataIn_1_valid_109;
  reg                 _zz_io_dataIn_1_valid_110;
  reg                 _zz_io_dataIn_1_valid_111;
  reg                 _zz_io_dataIn_1_valid_112;
  reg                 _zz_io_dataIn_1_valid_113;
  reg                 _zz_io_dataIn_1_valid_114;
  reg                 _zz_io_dataIn_1_valid_115;
  reg                 _zz_io_dataIn_1_valid_116;
  reg                 _zz_io_dataIn_1_valid_117;
  reg                 _zz_io_dataIn_1_valid_118;
  reg                 _zz_io_dataIn_1_valid_119;
  reg                 _zz_io_dataIn_1_valid_120;
  reg                 _zz_io_dataIn_1_valid_121;
  reg                 _zz_io_dataIn_1_valid_122;
  reg                 _zz_io_dataIn_1_valid_123;
  reg                 _zz_io_dataIn_1_valid_124;
  reg                 _zz_io_dataIn_1_valid_125;
  reg                 _zz_io_dataIn_1_valid_126;
  reg                 _zz_io_dataIn_1_valid_127;
  reg                 _zz_io_dataIn_1_valid_128;
  reg                 _zz_io_dataIn_1_valid_129;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_X;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_Y;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_Z;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_T;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_30;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_31;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_32;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_33;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_34;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_35;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_36;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_37;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_38;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_39;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_40;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_41;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_42;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_43;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_44;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_45;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_46;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_47;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_48;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_49;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_50;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_51;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_52;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_53;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_54;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_55;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_56;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_57;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_58;
  reg        [15:0]   _zz_io_dataIn_1_payload_address_59;
  wire                when_Pippenger_l207;
  reg                 _zz_io_dataIn_1_valid_130;
  reg                 _zz_io_dataIn_1_valid_131;
  reg                 _zz_io_dataIn_1_valid_132;
  reg                 _zz_io_dataIn_1_valid_133;
  reg                 _zz_io_dataIn_1_valid_134;
  reg                 _zz_io_dataIn_1_valid_135;
  reg                 _zz_io_dataIn_1_valid_136;
  reg                 _zz_io_dataIn_1_valid_137;
  reg                 _zz_io_dataIn_1_valid_138;
  reg                 _zz_io_dataIn_1_valid_139;
  reg                 _zz_io_dataIn_1_valid_140;
  reg                 _zz_io_dataIn_1_valid_141;
  reg                 _zz_io_dataIn_1_valid_142;
  reg                 _zz_io_dataIn_1_valid_143;
  reg                 _zz_io_dataIn_1_valid_144;
  reg                 _zz_io_dataIn_1_valid_145;
  reg                 _zz_io_dataIn_1_valid_146;
  reg                 _zz_io_dataIn_1_valid_147;
  reg                 _zz_io_dataIn_1_valid_148;
  reg                 _zz_io_dataIn_1_valid_149;
  reg                 _zz_io_dataIn_1_valid_150;
  reg                 _zz_io_dataIn_1_valid_151;
  reg                 _zz_io_dataIn_1_valid_152;
  reg                 _zz_io_dataIn_1_valid_153;
  reg                 _zz_io_dataIn_1_valid_154;
  reg                 _zz_io_dataIn_1_valid_155;
  reg                 _zz_io_dataIn_1_valid_156;
  reg                 _zz_io_dataIn_1_valid_157;
  reg                 _zz_io_dataIn_1_valid_158;
  reg                 _zz_io_dataIn_1_valid_159;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_X_1;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_Y_1;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_Z_1;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_T_1;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_60;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_61;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_62;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_63;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_64;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_65;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_66;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_67;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_68;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_69;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_70;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_71;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_72;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_73;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_74;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_75;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_76;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_77;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_78;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_79;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_80;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_81;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_82;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_83;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_84;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_85;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_86;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_87;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_88;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_89;
  reg                 _zz_io_dataIn_1_valid_160;
  reg                 _zz_io_dataIn_1_valid_161;
  reg                 _zz_io_dataIn_1_valid_162;
  reg                 _zz_io_dataIn_1_valid_163;
  reg                 _zz_io_dataIn_1_valid_164;
  reg                 _zz_io_dataIn_1_valid_165;
  reg                 _zz_io_dataIn_1_valid_166;
  reg                 _zz_io_dataIn_1_valid_167;
  reg                 _zz_io_dataIn_1_valid_168;
  reg                 _zz_io_dataIn_1_valid_169;
  reg                 _zz_io_dataIn_1_valid_170;
  reg                 _zz_io_dataIn_1_valid_171;
  reg                 _zz_io_dataIn_1_valid_172;
  reg                 _zz_io_dataIn_1_valid_173;
  reg                 _zz_io_dataIn_1_valid_174;
  reg                 _zz_io_dataIn_1_valid_175;
  reg                 _zz_io_dataIn_1_valid_176;
  reg                 _zz_io_dataIn_1_valid_177;
  reg                 _zz_io_dataIn_1_valid_178;
  reg                 _zz_io_dataIn_1_valid_179;
  reg                 _zz_io_dataIn_1_valid_180;
  reg                 _zz_io_dataIn_1_valid_181;
  reg                 _zz_io_dataIn_1_valid_182;
  reg                 _zz_io_dataIn_1_valid_183;
  reg                 _zz_io_dataIn_1_valid_184;
  reg                 _zz_io_dataIn_1_valid_185;
  reg                 _zz_io_dataIn_1_valid_186;
  reg                 _zz_io_dataIn_1_valid_187;
  reg                 _zz_io_dataIn_1_valid_188;
  reg                 _zz_io_dataIn_1_valid_189;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_X_1;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_1;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_1;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_T_1;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_90;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_91;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_92;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_93;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_94;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_95;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_96;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_97;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_98;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_99;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_100;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_101;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_102;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_103;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_104;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_105;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_106;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_107;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_108;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_109;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_110;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_111;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_112;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_113;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_114;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_115;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_116;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_117;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_118;
  reg        [3:0]    _zz_io_dataIn_1_payload_address_119;
  wire                when_Pippenger_l249;
  reg                 _zz_io_dataIn_1_valid_190;
  reg                 _zz_io_dataIn_1_valid_191;
  reg                 _zz_io_dataIn_1_valid_192;
  reg                 _zz_io_dataIn_1_valid_193;
  reg                 _zz_io_dataIn_1_valid_194;
  reg                 _zz_io_dataIn_1_valid_195;
  reg                 _zz_io_dataIn_1_valid_196;
  reg                 _zz_io_dataIn_1_valid_197;
  reg                 _zz_io_dataIn_1_valid_198;
  reg                 _zz_io_dataIn_1_valid_199;
  reg                 _zz_io_dataIn_1_valid_200;
  reg                 _zz_io_dataIn_1_valid_201;
  reg                 _zz_io_dataIn_1_valid_202;
  reg                 _zz_io_dataIn_1_valid_203;
  reg                 _zz_io_dataIn_1_valid_204;
  reg                 _zz_io_dataIn_1_valid_205;
  reg                 _zz_io_dataIn_1_valid_206;
  reg                 _zz_io_dataIn_1_valid_207;
  reg                 _zz_io_dataIn_1_valid_208;
  reg                 _zz_io_dataIn_1_valid_209;
  reg                 _zz_io_dataIn_1_valid_210;
  reg                 _zz_io_dataIn_1_valid_211;
  reg                 _zz_io_dataIn_1_valid_212;
  reg                 _zz_io_dataIn_1_valid_213;
  reg                 _zz_io_dataIn_1_valid_214;
  reg                 _zz_io_dataIn_1_valid_215;
  reg                 _zz_io_dataIn_1_valid_216;
  reg                 _zz_io_dataIn_1_valid_217;
  reg                 _zz_io_dataIn_1_valid_218;
  reg                 _zz_io_dataIn_1_valid_219;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_X_2;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_2;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_2;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_T_2;
  reg                 _zz_io_dataIn_1_valid_220;
  reg                 _zz_io_dataIn_1_valid_221;
  reg                 _zz_io_dataIn_1_valid_222;
  reg                 _zz_io_dataIn_1_valid_223;
  reg                 _zz_io_dataIn_1_valid_224;
  reg                 _zz_io_dataIn_1_valid_225;
  reg                 _zz_io_dataIn_1_valid_226;
  reg                 _zz_io_dataIn_1_valid_227;
  reg                 _zz_io_dataIn_1_valid_228;
  reg                 _zz_io_dataIn_1_valid_229;
  reg                 _zz_io_dataIn_1_valid_230;
  reg                 _zz_io_dataIn_1_valid_231;
  reg                 _zz_io_dataIn_1_valid_232;
  reg                 _zz_io_dataIn_1_valid_233;
  reg                 _zz_io_dataIn_1_valid_234;
  reg                 _zz_io_dataIn_1_valid_235;
  reg                 _zz_io_dataIn_1_valid_236;
  reg                 _zz_io_dataIn_1_valid_237;
  reg                 _zz_io_dataIn_1_valid_238;
  reg                 _zz_io_dataIn_1_valid_239;
  reg                 _zz_io_dataIn_1_valid_240;
  reg                 _zz_io_dataIn_1_valid_241;
  reg                 _zz_io_dataIn_1_valid_242;
  reg                 _zz_io_dataIn_1_valid_243;
  reg                 _zz_io_dataIn_1_valid_244;
  reg                 _zz_io_dataIn_1_valid_245;
  reg                 _zz_io_dataIn_1_valid_246;
  reg                 _zz_io_dataIn_1_valid_247;
  reg                 _zz_io_dataIn_1_valid_248;
  reg                 _zz_io_dataIn_1_valid_249;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_X_3;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_3;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_3;
  reg        [376:0]  pippenger_1_dataRam_1_1_io_rData_1_regNext_T_3;
  wire                when_Pippenger_l306;
  wire                when_Pippenger_l319;
  `ifndef SYNTHESIS
  reg [87:0] fsm_stateReg_string;
  reg [87:0] fsm_stateNext_string;
  `endif


  assign _zz_dataInBuffer_dataReg_fragment_K = (dataInBuffer_dataReg_fragment_K >>> 26);
  assign _zz_flushing_flushCnt_valueNext_1 = flushing_flushCnt_willIncrement;
  assign _zz_flushing_flushCnt_valueNext = {15'd0, _zz_flushing_flushCnt_valueNext_1};
  assign _zz_stage1_NCnt_valueNext_1 = stage1_NCnt_willIncrement;
  assign _zz_stage1_NCnt_valueNext = {31'd0, _zz_stage1_NCnt_valueNext_1};
  assign _zz_stage1_GCnt_valueNext_1 = stage1_GCnt_willIncrement;
  assign _zz_stage1_GCnt_valueNext = {3'd0, _zz_stage1_GCnt_valueNext_1};
  assign _zz_stage1_emptyCnt_valueNext_1 = stage1_emptyCnt_willIncrement;
  assign _zz_stage1_emptyCnt_valueNext = {8'd0, _zz_stage1_emptyCnt_valueNext_1};
  assign _zz_stage1_inputBarrelID_0_2 = {1'b0,stage1_needAdd1_0};
  assign _zz_stage1_inputBarrelID_0_1 = {12'd0, _zz_stage1_inputBarrelID_0_2};
  assign _zz_stage1_inputBarrelID_1_1 = {1'b0,(|stage1_inputBarrelID_0[13 : 12])};
  assign _zz_stage1_inputBarrelID_1 = {12'd0, _zz_stage1_inputBarrelID_1_1};
  assign _zz__zz_stage1_inputBarrelIDAbs_0 = stage1_inputBarrelID_0[12:0];
  assign _zz_stage1_inputBarrelIDAbs_0_1 = (_zz_stage1_inputBarrelIDAbs_0_2 + _zz_stage1_inputBarrelIDAbs_0_4);
  assign _zz_stage1_inputBarrelIDAbs_0_2 = (_zz_stage1_inputBarrelIDAbs_0[12] ? _zz_stage1_inputBarrelIDAbs_0_3 : _zz_stage1_inputBarrelIDAbs_0);
  assign _zz_stage1_inputBarrelIDAbs_0_3 = (~ _zz_stage1_inputBarrelIDAbs_0);
  assign _zz_stage1_inputBarrelIDAbs_0_5 = _zz_stage1_inputBarrelIDAbs_0[12];
  assign _zz_stage1_inputBarrelIDAbs_0_4 = {12'd0, _zz_stage1_inputBarrelIDAbs_0_5};
  assign _zz__zz_stage1_inputBarrelIDAbs_1 = stage1_inputBarrelID_1[12:0];
  assign _zz_stage1_inputBarrelIDAbs_1_1 = (_zz_stage1_inputBarrelIDAbs_1_2 + _zz_stage1_inputBarrelIDAbs_1_4);
  assign _zz_stage1_inputBarrelIDAbs_1_2 = (_zz_stage1_inputBarrelIDAbs_1[12] ? _zz_stage1_inputBarrelIDAbs_1_3 : _zz_stage1_inputBarrelIDAbs_1);
  assign _zz_stage1_inputBarrelIDAbs_1_3 = (~ _zz_stage1_inputBarrelIDAbs_1);
  assign _zz_stage1_inputBarrelIDAbs_1_5 = _zz_stage1_inputBarrelIDAbs_1[12];
  assign _zz_stage1_inputBarrelIDAbs_1_4 = {12'd0, _zz_stage1_inputBarrelIDAbs_1_5};
  assign _zz__zz_stage1_inputValid_0 = stage1_inputBarrelID_0[12:0];
  assign _zz__zz_stage1_inputValid_1 = stage1_inputBarrelID_1[12:0];
  assign _zz_stage2_wCnt_valueNext_1 = stage2_wCnt_willDecrement;
  assign _zz_stage2_wCnt_valueNext = {11'd0, _zz_stage2_wCnt_valueNext_1};
  assign _zz_stage2_GCnt_valueNext_1 = stage2_GCnt_willIncrement;
  assign _zz_stage2_GCnt_valueNext = {3'd0, _zz_stage2_GCnt_valueNext_1};
  assign _zz_stage2_calCnt_valueNext_1 = stage2_calCnt_willDecrement;
  assign _zz_stage2_calCnt_valueNext = {1'd0, _zz_stage2_calCnt_valueNext_1};
  assign _zz_stage2_waitCnt_valueNext_1 = stage2_waitCnt_willIncrement;
  assign _zz_stage2_waitCnt_valueNext = {8'd0, _zz_stage2_waitCnt_valueNext_1};
  assign _zz_stage3_GCnt_valueNext_1 = stage3_GCnt_willDecrement;
  assign _zz_stage3_GCnt_valueNext = {3'd0, _zz_stage3_GCnt_valueNext_1};
  assign _zz_stage3_doubleCnt_valueNext_1 = stage3_doubleCnt_willIncrement;
  assign _zz_stage3_doubleCnt_valueNext = {4'd0, _zz_stage3_doubleCnt_valueNext_1};
  assign _zz_stage3_doubleWaitCnt_valueNext_1 = stage3_doubleWaitCnt_willIncrement;
  assign _zz_stage3_doubleWaitCnt_valueNext = {8'd0, _zz_stage3_doubleWaitCnt_valueNext_1};
  assign _zz_stage3_addWaitCnt_valueNext_1 = stage3_addWaitCnt_willIncrement;
  assign _zz_stage3_addWaitCnt_valueNext = {8'd0, _zz_stage3_addWaitCnt_valueNext_1};
  assign _zz_stage3Final_doubleCnt_valueNext_1 = stage3Final_doubleCnt_willIncrement;
  assign _zz_stage3Final_doubleCnt_valueNext = {3'd0, _zz_stage3Final_doubleCnt_valueNext_1};
  assign _zz_stage3Final_doubleWaitCnt_valueNext_1 = stage3Final_doubleWaitCnt_willIncrement;
  assign _zz_stage3Final_doubleWaitCnt_valueNext = {8'd0, _zz_stage3Final_doubleWaitCnt_valueNext_1};
  assign _zz_stage3Final_addWaitCnt_valueNext_1 = stage3Final_addWaitCnt_willIncrement;
  assign _zz_stage3Final_addWaitCnt_valueNext = {8'd0, _zz_stage3Final_addWaitCnt_valueNext_1};
  assign _zz_io_address_0_1 = (stage2_wCnt_value + _zz_io_address_0_2);
  assign _zz_io_address_0 = _zz_io_address_0_1;
  assign _zz_io_address_0_2 = {10'd0, stage2_calCnt_value};
  assign _zz_io_address_1_1 = (stage2_wCnt_value + _zz_io_address_1_2);
  assign _zz_io_address_1 = _zz_io_address_1_1;
  assign _zz_io_address_1_2 = {10'd0, stage2_calCnt_value};
  assign _zz__zz_io_dataIn_1_payload_address_1 = (stage2_wCnt_value + _zz__zz_io_dataIn_1_payload_address_2);
  assign _zz__zz_io_dataIn_1_payload_address = _zz__zz_io_dataIn_1_payload_address_1;
  assign _zz__zz_io_dataIn_1_payload_address_2 = {10'd0, stage2_calCnt_value};
  assign _zz_io_address_0_4 = (stage2_wCnt_value + _zz_io_address_0_5);
  assign _zz_io_address_0_3 = _zz_io_address_0_4;
  assign _zz_io_address_0_5 = {10'd0, stage2_calCnt_value};
  assign _zz_io_address_1_4 = (stage2_wCnt_value + _zz_io_address_1_5);
  assign _zz_io_address_1_3 = _zz_io_address_1_4;
  assign _zz_io_address_1_5 = {10'd0, stage2_calCnt_value};
  assign _zz__zz_io_dataIn_1_payload_address_30_1 = (stage2_wCnt_value + _zz__zz_io_dataIn_1_payload_address_30_2);
  assign _zz__zz_io_dataIn_1_payload_address_30 = _zz__zz_io_dataIn_1_payload_address_30_1;
  assign _zz__zz_io_dataIn_1_payload_address_30_2 = {10'd0, stage2_calCnt_value};
  assign _zz_io_address_1_6 = (stage3_GCnt_value - _zz_io_address_1_7);
  assign _zz_io_address_1_8 = stage3_addWaitCnt_value[0];
  assign _zz_io_address_1_7 = {3'd0, _zz_io_address_1_8};
  assign _zz__zz_io_dataIn_1_payload_address_60_1 = stage3_addWaitCnt_value[0];
  assign _zz__zz_io_dataIn_1_payload_address_60 = {3'd0, _zz__zz_io_dataIn_1_payload_address_60_1};
  assign _zz_io_address_1_9 = (stage3_GCnt_value - _zz_io_address_1_10);
  assign _zz_io_address_1_11 = stage3_addWaitCnt_value[0];
  assign _zz_io_address_1_10 = {3'd0, _zz_io_address_1_11};
  assign _zz__zz_io_dataIn_1_payload_address_90_1 = stage3_addWaitCnt_value[0];
  assign _zz__zz_io_dataIn_1_payload_address_90 = {3'd0, _zz__zz_io_dataIn_1_payload_address_90_1};
  StateRam stateRam_0 (
    .io_we_0      (stateRam_0_io_we_0           ), //i
    .io_we_1      (stateRam_0_io_we_1           ), //i
    .io_address_0 (stateRam_0_io_address_0[15:0]), //i
    .io_address_1 (stateRam_0_io_address_1[15:0]), //i
    .io_state_0   (stateRam_0_io_state_0        ), //o
    .io_state_1   (stateRam_0_io_state_1        ), //o
    .io_flush     (stateRam_0_io_flush          ), //i
    .io_flushCnt  (stateRam_0_io_flushCnt[15:0] ), //i
    .clk          (clk                          ), //i
    .resetn       (resetn                       )  //i
  );
  StateRam stateRam_1_1 (
    .io_we_0      (stateRam_1_1_io_we_0           ), //i
    .io_we_1      (stateRam_1_1_io_we_1           ), //i
    .io_address_0 (stateRam_1_1_io_address_0[15:0]), //i
    .io_address_1 (stateRam_1_1_io_address_1[15:0]), //i
    .io_state_0   (stateRam_1_1_io_state_0        ), //o
    .io_state_1   (stateRam_1_1_io_state_1        ), //o
    .io_flush     (stateRam_1_1_io_flush          ), //i
    .io_flushCnt  (stateRam_1_1_io_flushCnt[15:0] ), //i
    .clk          (clk                            ), //i
    .resetn       (resetn                         )  //i
  );
  DataRam dataRam_0 (
    .io_we_0      (dataRam_0_io_we_0            ), //i
    .io_we_1      (dataRam_0_io_we_1            ), //i
    .io_address_0 (dataRam_0_io_address_0[15:0] ), //i
    .io_address_1 (dataRam_0_io_address_1[15:0] ), //i
    .io_wData_0_X (dataRam_0_io_wData_0_X[376:0]), //i
    .io_wData_0_Y (dataRam_0_io_wData_0_Y[376:0]), //i
    .io_wData_0_Z (dataRam_0_io_wData_0_Z[376:0]), //i
    .io_wData_0_T (dataRam_0_io_wData_0_T[376:0]), //i
    .io_wData_1_X (dataRam_0_io_wData_1_X[376:0]), //i
    .io_wData_1_Y (dataRam_0_io_wData_1_Y[376:0]), //i
    .io_wData_1_Z (dataRam_0_io_wData_1_Z[376:0]), //i
    .io_wData_1_T (dataRam_0_io_wData_1_T[376:0]), //i
    .io_state_0   (1'b1                         ), //i
    .io_state_1   (dataRam_0_io_state_1         ), //i
    .io_rData_0_X (dataRam_0_io_rData_0_X[376:0]), //o
    .io_rData_0_Y (dataRam_0_io_rData_0_Y[376:0]), //o
    .io_rData_0_Z (dataRam_0_io_rData_0_Z[376:0]), //o
    .io_rData_0_T (dataRam_0_io_rData_0_T[376:0]), //o
    .io_rData_1_X (dataRam_0_io_rData_1_X[376:0]), //o
    .io_rData_1_Y (dataRam_0_io_rData_1_Y[376:0]), //o
    .io_rData_1_Z (dataRam_0_io_rData_1_Z[376:0]), //o
    .io_rData_1_T (dataRam_0_io_rData_1_T[376:0]), //o
    .io_pInit_X   (io_pInit_X[376:0]            ), //i
    .io_pInit_Y   (io_pInit_Y[376:0]            ), //i
    .io_pInit_Z   (io_pInit_Z[376:0]            ), //i
    .io_pInit_T   (io_pInit_T[376:0]            ), //i
    .clk          (clk                          ), //i
    .resetn       (resetn                       )  //i
  );
  DataRam dataRam_1_1 (
    .io_we_0      (dataRam_1_1_io_we_0            ), //i
    .io_we_1      (dataRam_1_1_io_we_1            ), //i
    .io_address_0 (dataRam_1_1_io_address_0[15:0] ), //i
    .io_address_1 (dataRam_1_1_io_address_1[15:0] ), //i
    .io_wData_0_X (dataRam_1_1_io_wData_0_X[376:0]), //i
    .io_wData_0_Y (dataRam_1_1_io_wData_0_Y[376:0]), //i
    .io_wData_0_Z (dataRam_1_1_io_wData_0_Z[376:0]), //i
    .io_wData_0_T (dataRam_1_1_io_wData_0_T[376:0]), //i
    .io_wData_1_X (dataRam_1_1_io_wData_1_X[376:0]), //i
    .io_wData_1_Y (dataRam_1_1_io_wData_1_Y[376:0]), //i
    .io_wData_1_Z (dataRam_1_1_io_wData_1_Z[376:0]), //i
    .io_wData_1_T (dataRam_1_1_io_wData_1_T[376:0]), //i
    .io_state_0   (1'b1                           ), //i
    .io_state_1   (dataRam_1_1_io_state_1         ), //i
    .io_rData_0_X (dataRam_1_1_io_rData_0_X[376:0]), //o
    .io_rData_0_Y (dataRam_1_1_io_rData_0_Y[376:0]), //o
    .io_rData_0_Z (dataRam_1_1_io_rData_0_Z[376:0]), //o
    .io_rData_0_T (dataRam_1_1_io_rData_0_T[376:0]), //o
    .io_rData_1_X (dataRam_1_1_io_rData_1_X[376:0]), //o
    .io_rData_1_Y (dataRam_1_1_io_rData_1_Y[376:0]), //o
    .io_rData_1_Z (dataRam_1_1_io_rData_1_Z[376:0]), //o
    .io_rData_1_T (dataRam_1_1_io_rData_1_T[376:0]), //o
    .io_pInit_X   (io_pInit_X[376:0]              ), //i
    .io_pInit_Y   (io_pInit_Y[376:0]              ), //i
    .io_pInit_Z   (io_pInit_Z[376:0]              ), //i
    .io_pInit_T   (io_pInit_T[376:0]              ), //i
    .clk          (clk                            ), //i
    .resetn       (resetn                         )  //i
  );
  DWSRFIFO fifo_0 (
    .io_dataIn_0_valid           (fifo_0_io_dataIn_0_valid                ), //i
    .io_dataIn_0_payload_a_X     (fifo_0_io_dataIn_0_payload_a_X[376:0]   ), //i
    .io_dataIn_0_payload_a_Y     (fifo_0_io_dataIn_0_payload_a_Y[376:0]   ), //i
    .io_dataIn_0_payload_a_Z     (fifo_0_io_dataIn_0_payload_a_Z[376:0]   ), //i
    .io_dataIn_0_payload_a_T     (fifo_0_io_dataIn_0_payload_a_T[376:0]   ), //i
    .io_dataIn_0_payload_b_X     (fifo_0_io_dataIn_0_payload_b_X[376:0]   ), //i
    .io_dataIn_0_payload_b_Y     (fifo_0_io_dataIn_0_payload_b_Y[376:0]   ), //i
    .io_dataIn_0_payload_b_Z     (fifo_0_io_dataIn_0_payload_b_Z[376:0]   ), //i
    .io_dataIn_0_payload_b_T     (fifo_0_io_dataIn_0_payload_b_T[376:0]   ), //i
    .io_dataIn_0_payload_address (fifo_0_io_dataIn_0_payload_address[15:0]), //i
    .io_dataIn_1_valid           (fifo_0_io_dataIn_1_valid                ), //i
    .io_dataIn_1_payload_a_X     (fifo_0_io_dataIn_1_payload_a_X[376:0]   ), //i
    .io_dataIn_1_payload_a_Y     (fifo_0_io_dataIn_1_payload_a_Y[376:0]   ), //i
    .io_dataIn_1_payload_a_Z     (fifo_0_io_dataIn_1_payload_a_Z[376:0]   ), //i
    .io_dataIn_1_payload_a_T     (fifo_0_io_dataIn_1_payload_a_T[376:0]   ), //i
    .io_dataIn_1_payload_b_X     (fifo_0_io_dataIn_1_payload_b_X[376:0]   ), //i
    .io_dataIn_1_payload_b_Y     (fifo_0_io_dataIn_1_payload_b_Y[376:0]   ), //i
    .io_dataIn_1_payload_b_Z     (fifo_0_io_dataIn_1_payload_b_Z[376:0]   ), //i
    .io_dataIn_1_payload_b_T     (fifo_0_io_dataIn_1_payload_b_T[376:0]   ), //i
    .io_dataIn_1_payload_address (fifo_0_io_dataIn_1_payload_address[15:0]), //i
    .io_dataOut_valid            (fifo_0_io_dataOut_valid                 ), //o
    .io_dataOut_payload_a_X      (fifo_0_io_dataOut_payload_a_X[376:0]    ), //o
    .io_dataOut_payload_a_Y      (fifo_0_io_dataOut_payload_a_Y[376:0]    ), //o
    .io_dataOut_payload_a_Z      (fifo_0_io_dataOut_payload_a_Z[376:0]    ), //o
    .io_dataOut_payload_a_T      (fifo_0_io_dataOut_payload_a_T[376:0]    ), //o
    .io_dataOut_payload_b_X      (fifo_0_io_dataOut_payload_b_X[376:0]    ), //o
    .io_dataOut_payload_b_Y      (fifo_0_io_dataOut_payload_b_Y[376:0]    ), //o
    .io_dataOut_payload_b_Z      (fifo_0_io_dataOut_payload_b_Z[376:0]    ), //o
    .io_dataOut_payload_b_T      (fifo_0_io_dataOut_payload_b_T[376:0]    ), //o
    .io_dataOut_payload_address  (fifo_0_io_dataOut_payload_address[15:0] ), //o
    .clk                         (clk                                     ), //i
    .resetn                      (resetn                                  )  //i
  );
  DWSRFIFO fifo_1 (
    .io_dataIn_0_valid           (fifo_1_io_dataIn_0_valid                ), //i
    .io_dataIn_0_payload_a_X     (fifo_1_io_dataIn_0_payload_a_X[376:0]   ), //i
    .io_dataIn_0_payload_a_Y     (fifo_1_io_dataIn_0_payload_a_Y[376:0]   ), //i
    .io_dataIn_0_payload_a_Z     (fifo_1_io_dataIn_0_payload_a_Z[376:0]   ), //i
    .io_dataIn_0_payload_a_T     (fifo_1_io_dataIn_0_payload_a_T[376:0]   ), //i
    .io_dataIn_0_payload_b_X     (fifo_1_io_dataIn_0_payload_b_X[376:0]   ), //i
    .io_dataIn_0_payload_b_Y     (fifo_1_io_dataIn_0_payload_b_Y[376:0]   ), //i
    .io_dataIn_0_payload_b_Z     (fifo_1_io_dataIn_0_payload_b_Z[376:0]   ), //i
    .io_dataIn_0_payload_b_T     (fifo_1_io_dataIn_0_payload_b_T[376:0]   ), //i
    .io_dataIn_0_payload_address (fifo_1_io_dataIn_0_payload_address[15:0]), //i
    .io_dataIn_1_valid           (fifo_1_io_dataIn_1_valid                ), //i
    .io_dataIn_1_payload_a_X     (fifo_1_io_dataIn_1_payload_a_X[376:0]   ), //i
    .io_dataIn_1_payload_a_Y     (fifo_1_io_dataIn_1_payload_a_Y[376:0]   ), //i
    .io_dataIn_1_payload_a_Z     (fifo_1_io_dataIn_1_payload_a_Z[376:0]   ), //i
    .io_dataIn_1_payload_a_T     (fifo_1_io_dataIn_1_payload_a_T[376:0]   ), //i
    .io_dataIn_1_payload_b_X     (fifo_1_io_dataIn_1_payload_b_X[376:0]   ), //i
    .io_dataIn_1_payload_b_Y     (fifo_1_io_dataIn_1_payload_b_Y[376:0]   ), //i
    .io_dataIn_1_payload_b_Z     (fifo_1_io_dataIn_1_payload_b_Z[376:0]   ), //i
    .io_dataIn_1_payload_b_T     (fifo_1_io_dataIn_1_payload_b_T[376:0]   ), //i
    .io_dataIn_1_payload_address (fifo_1_io_dataIn_1_payload_address[15:0]), //i
    .io_dataOut_valid            (fifo_1_io_dataOut_valid                 ), //o
    .io_dataOut_payload_a_X      (fifo_1_io_dataOut_payload_a_X[376:0]    ), //o
    .io_dataOut_payload_a_Y      (fifo_1_io_dataOut_payload_a_Y[376:0]    ), //o
    .io_dataOut_payload_a_Z      (fifo_1_io_dataOut_payload_a_Z[376:0]    ), //o
    .io_dataOut_payload_a_T      (fifo_1_io_dataOut_payload_a_T[376:0]    ), //o
    .io_dataOut_payload_b_X      (fifo_1_io_dataOut_payload_b_X[376:0]    ), //o
    .io_dataOut_payload_b_Y      (fifo_1_io_dataOut_payload_b_Y[376:0]    ), //o
    .io_dataOut_payload_b_Z      (fifo_1_io_dataOut_payload_b_Z[376:0]    ), //o
    .io_dataOut_payload_b_T      (fifo_1_io_dataOut_payload_b_T[376:0]    ), //o
    .io_dataOut_payload_address  (fifo_1_io_dataOut_payload_address[15:0] ), //o
    .clk                         (clk                                     ), //i
    .resetn                      (resetn                                  )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_flushing : fsm_stateReg_string = "flushing   ";
      fsm_enumDef_stage1 : fsm_stateReg_string = "stage1     ";
      fsm_enumDef_stage2 : fsm_stateReg_string = "stage2     ";
      fsm_enumDef_stage3 : fsm_stateReg_string = "stage3     ";
      fsm_enumDef_stage3Final : fsm_stateReg_string = "stage3Final";
      default : fsm_stateReg_string = "???????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_flushing : fsm_stateNext_string = "flushing   ";
      fsm_enumDef_stage1 : fsm_stateNext_string = "stage1     ";
      fsm_enumDef_stage2 : fsm_stateNext_string = "stage2     ";
      fsm_enumDef_stage3 : fsm_stateNext_string = "stage3     ";
      fsm_enumDef_stage3Final : fsm_stateNext_string = "stage3Final";
      default : fsm_stateNext_string = "???????????";
    endcase
  end
  `endif

  assign dataInBuffer_bufferOut_valid = dataInBuffer_validReg;
  assign dataInBuffer_bufferOut_payload_last = dataInBuffer_dataReg_last;
  assign dataInBuffer_bufferOut_payload_fragment_P_X = dataInBuffer_dataReg_fragment_P_X;
  assign dataInBuffer_bufferOut_payload_fragment_P_Y = dataInBuffer_dataReg_fragment_P_Y;
  assign dataInBuffer_bufferOut_payload_fragment_P_Z = dataInBuffer_dataReg_fragment_P_Z;
  assign dataInBuffer_bufferOut_payload_fragment_P_T = dataInBuffer_dataReg_fragment_P_T;
  assign dataInBuffer_bufferOut_payload_fragment_K = dataInBuffer_dataReg_fragment_K;
  assign io_dataIn_ready = ((! dataInBuffer_validReg) || dataInBuffer_bufferOut_ready);
  always @(*) begin
    dataInBuffer_bufferOut_ready = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          if(dataInBuffer_bufferOut_valid) begin
            if(stage1_GCnt_willOverflowIfInc) begin
              dataInBuffer_bufferOut_ready = 1'b1;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataInBuffer_shift = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          dataInBuffer_shift = 1'b1;
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_we_0 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_0_io_we_0 = shiftRegs_validOut_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_we_1 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_0_io_we_1 = stage1_inputValid_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_1_1_io_we_0 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_1_1_io_we_0 = shiftRegs_validOut_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_1_1_io_we_1 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_1_1_io_we_1 = stage1_inputValid_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_address_0 = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_0_io_address_0 = shiftRegs_addressOut_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_0_io_address_0 = {stage2_GCnt_value,_zz_io_address_0};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_address_1 = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_0_io_address_1 = stage1_inputAddress_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_1_1_io_address_0 = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_1_1_io_address_0 = shiftRegs_addressOut_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_1_1_io_address_0 = {stage2_GCnt_value,_zz_io_address_0_3};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_1_1_io_address_1 = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_1_1_io_address_1 = stage1_inputAddress_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_flush = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_0_io_flush = stage2_calCnt_willUnderflowIfDec;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
        stateRam_0_io_flush = 1'b1;
      end
    endcase
  end

  always @(*) begin
    stateRam_1_1_io_flush = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_1_1_io_flush = stage2_calCnt_willUnderflowIfDec;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
        stateRam_1_1_io_flush = 1'b1;
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_flushCnt = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_0_io_flushCnt = {stage2_GCnt_value,stage2_wCnt_value};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
        stateRam_0_io_flushCnt = flushing_flushCnt_value;
      end
    endcase
  end

  always @(*) begin
    stateRam_1_1_io_flushCnt = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_1_1_io_flushCnt = {stage2_GCnt_value,stage2_wCnt_value};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
        stateRam_1_1_io_flushCnt = flushing_flushCnt_value;
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_we_0 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_we_0 = ((! stateRam_0_io_state_0) && shiftRegs_validOutFull_0);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_we_0 = shiftRegs_validOutFull_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_we_0 = shiftRegs_validOutFull_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_we_1 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_we_1 = ((! stateRam_0_io_state_1) && stage1_inputValid_0_delay_5);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_we_0 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_we_0 = ((! stateRam_1_1_io_state_0) && shiftRegs_validOutFull_1);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_1_1_io_we_0 = shiftRegs_validOutFull_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_1_1_io_we_0 = shiftRegs_validOutFull_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        dataRam_1_1_io_we_0 = shiftRegs_validOutFull_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_we_1 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_we_1 = ((! stateRam_1_1_io_state_1) && stage1_inputValid_1_delay_5);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_address_0 = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_address_0 = shiftRegs_addressOutFull_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_address_0 = shiftRegs_addressOutFull_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_address_0 = shiftRegs_addressOutFull_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_address_1 = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_address_1 = stage1_inputAddress_0_delay_5;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_address_1 = {stage2_GCnt_value,_zz_io_address_1};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_address_1 = {_zz_io_address_1_6,12'h001};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        dataRam_0_io_address_1 = 16'h0001;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_address_0 = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_address_0 = shiftRegs_addressOutFull_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_1_1_io_address_0 = shiftRegs_addressOutFull_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_1_1_io_address_0 = shiftRegs_addressOutFull_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        dataRam_1_1_io_address_0 = shiftRegs_addressOutFull_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_address_1 = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_address_1 = stage1_inputAddress_1_delay_5;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_1_1_io_address_1 = {stage2_GCnt_value,_zz_io_address_1_3};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_1_1_io_address_1 = {_zz_io_address_1_9,12'h001};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        dataRam_1_1_io_address_1 = 16'h0001;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_0_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_0_X = pAddPort_0_s_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_wData_0_X = pAddPort_0_s_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_wData_0_X = pAddPort_0_s_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_0_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_0_Y = pAddPort_0_s_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_wData_0_Y = pAddPort_0_s_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_wData_0_Y = pAddPort_0_s_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_0_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_0_Z = pAddPort_0_s_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_wData_0_Z = pAddPort_0_s_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_wData_0_Z = pAddPort_0_s_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_0_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_0_T = pAddPort_0_s_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_wData_0_T = pAddPort_0_s_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_wData_0_T = pAddPort_0_s_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_1_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_1_X = stage1_inputData_0_delay_5_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_1_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_1_Y = stage1_inputData_0_delay_5_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_1_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_1_Z = stage1_inputData_0_delay_5_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_1_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_1_T = stage1_inputData_0_delay_5_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_wData_0_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_wData_0_X = pAddPort_1_s_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_1_1_io_wData_0_X = pAddPort_1_s_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_1_1_io_wData_0_X = pAddPort_1_s_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        dataRam_1_1_io_wData_0_X = pAddPort_1_s_X;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_wData_0_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_wData_0_Y = pAddPort_1_s_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_1_1_io_wData_0_Y = pAddPort_1_s_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_1_1_io_wData_0_Y = pAddPort_1_s_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        dataRam_1_1_io_wData_0_Y = pAddPort_1_s_Y;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_wData_0_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_wData_0_Z = pAddPort_1_s_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_1_1_io_wData_0_Z = pAddPort_1_s_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_1_1_io_wData_0_Z = pAddPort_1_s_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        dataRam_1_1_io_wData_0_Z = pAddPort_1_s_Z;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_wData_0_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_wData_0_T = pAddPort_1_s_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_1_1_io_wData_0_T = pAddPort_1_s_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_1_1_io_wData_0_T = pAddPort_1_s_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        dataRam_1_1_io_wData_0_T = pAddPort_1_s_T;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_wData_1_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_wData_1_X = stage1_inputData_1_delay_5_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_wData_1_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_wData_1_Y = stage1_inputData_1_delay_5_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_wData_1_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_wData_1_Z = stage1_inputData_1_delay_5_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_wData_1_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_1_1_io_wData_1_T = stage1_inputData_1_delay_5_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_state_1 = 1'b1;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_state_1 = _zz_io_state_1_38;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_1_1_io_state_1 = 1'b1;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_1_1_io_state_1 = _zz_io_state_1_77;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_valid = _zz_io_dataIn_0_valid_34;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_a_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_a_X = (_zz_io_dataIn_0_payload_a_X_34 ? stage1_inputData_0_delay_35_X : dataRam_0_io_rData_0_X);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_a_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_a_Y = (_zz_io_dataIn_0_payload_a_X_34 ? stage1_inputData_0_delay_35_Y : dataRam_0_io_rData_0_Y);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_a_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_a_Z = (_zz_io_dataIn_0_payload_a_X_34 ? stage1_inputData_0_delay_35_Z : dataRam_0_io_rData_0_Z);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_a_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_a_T = (_zz_io_dataIn_0_payload_a_X_34 ? stage1_inputData_0_delay_35_T : dataRam_0_io_rData_0_T);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_b_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_b_X = pAddPort_0_s_delay_30_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_b_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_b_Y = pAddPort_0_s_delay_30_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_b_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_b_Z = pAddPort_0_s_delay_30_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_b_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_b_T = pAddPort_0_s_delay_30_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_address = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_address = shiftRegs_addressOutFull_0_delay_30;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_valid = _zz_io_dataIn_1_valid_34;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_valid = _zz_io_dataIn_1_valid_99;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_valid = _zz_io_dataIn_1_valid_159;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_valid = _zz_io_dataIn_1_valid_219;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_a_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_a_X = dataRam_0_io_rData_1_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_a_X = dataRam_0_io_rData_1_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_a_X = dataRam_0_io_rData_1_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_payload_a_X = dataRam_0_io_rData_1_X;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_a_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_a_Y = dataRam_0_io_rData_1_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_a_Y = dataRam_0_io_rData_1_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_a_Y = dataRam_0_io_rData_1_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_payload_a_Y = dataRam_0_io_rData_1_Y;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_a_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_a_Z = dataRam_0_io_rData_1_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_a_Z = dataRam_0_io_rData_1_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_a_Z = dataRam_0_io_rData_1_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_payload_a_Z = dataRam_0_io_rData_1_Z;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_a_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_a_T = dataRam_0_io_rData_1_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_a_T = dataRam_0_io_rData_1_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_a_T = dataRam_0_io_rData_1_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_payload_a_T = dataRam_0_io_rData_1_T;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_b_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_b_X = stage1_inputData_0_delay_35_X_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_b_X = pippenger_1_dataRam_0_io_rData_1_regNext_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_b_X = pippenger_1_dataRam_0_io_rData_1_regNext_X_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_payload_b_X = pippenger_1_dataRam_1_1_io_rData_1_regNext_X_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_b_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_b_Y = stage1_inputData_0_delay_35_Y_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_b_Y = pippenger_1_dataRam_0_io_rData_1_regNext_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_b_Y = pippenger_1_dataRam_0_io_rData_1_regNext_Y_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_payload_b_Y = pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_b_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_b_Z = stage1_inputData_0_delay_35_Z_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_b_Z = pippenger_1_dataRam_0_io_rData_1_regNext_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_b_Z = pippenger_1_dataRam_0_io_rData_1_regNext_Z_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_payload_b_Z = pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_b_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_b_T = stage1_inputData_0_delay_35_T_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_b_T = pippenger_1_dataRam_0_io_rData_1_regNext_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_b_T = pippenger_1_dataRam_0_io_rData_1_regNext_T_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_0_io_dataIn_1_payload_b_T = pippenger_1_dataRam_1_1_io_rData_1_regNext_T_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_address = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_address = stage1_inputAddress_0_delay_35;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_address = _zz_io_dataIn_1_payload_address_29;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_address = {_zz_io_dataIn_1_payload_address_89,12'h001};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_valid = _zz_io_dataIn_0_valid_69;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_a_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_a_X = (_zz_io_dataIn_0_payload_a_X_69 ? stage1_inputData_1_delay_35_X : dataRam_1_1_io_rData_0_X);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_a_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_a_Y = (_zz_io_dataIn_0_payload_a_X_69 ? stage1_inputData_1_delay_35_Y : dataRam_1_1_io_rData_0_Y);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_a_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_a_Z = (_zz_io_dataIn_0_payload_a_X_69 ? stage1_inputData_1_delay_35_Z : dataRam_1_1_io_rData_0_Z);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_a_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_a_T = (_zz_io_dataIn_0_payload_a_X_69 ? stage1_inputData_1_delay_35_T : dataRam_1_1_io_rData_0_T);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_b_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_b_X = pAddPort_1_s_delay_30_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_b_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_b_Y = pAddPort_1_s_delay_30_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_b_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_b_Z = pAddPort_1_s_delay_30_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_b_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_b_T = pAddPort_1_s_delay_30_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_0_payload_address = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_0_payload_address = shiftRegs_addressOutFull_1_delay_30;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_valid = _zz_io_dataIn_1_valid_69;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_valid = _zz_io_dataIn_1_valid_129;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_valid = _zz_io_dataIn_1_valid_189;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_valid = _zz_io_dataIn_1_valid_249;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_a_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_a_X = dataRam_1_1_io_rData_1_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_a_X = dataRam_1_1_io_rData_1_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_a_X = dataRam_1_1_io_rData_1_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_a_X = dataRam_1_1_io_rData_1_X;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_a_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_a_Y = dataRam_1_1_io_rData_1_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_a_Y = dataRam_1_1_io_rData_1_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_a_Y = dataRam_1_1_io_rData_1_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_a_Y = dataRam_1_1_io_rData_1_Y;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_a_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_a_Z = dataRam_1_1_io_rData_1_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_a_Z = dataRam_1_1_io_rData_1_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_a_Z = dataRam_1_1_io_rData_1_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_a_Z = dataRam_1_1_io_rData_1_Z;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_a_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_a_T = dataRam_1_1_io_rData_1_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_a_T = dataRam_1_1_io_rData_1_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_a_T = dataRam_1_1_io_rData_1_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_a_T = dataRam_1_1_io_rData_1_T;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_b_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_b_X = stage1_inputData_1_delay_35_X_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_b_X = pippenger_1_dataRam_1_1_io_rData_1_regNext_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_b_X = pippenger_1_dataRam_1_1_io_rData_1_regNext_X_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_b_X = pippenger_1_dataRam_1_1_io_rData_1_regNext_X_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_b_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_b_Y = stage1_inputData_1_delay_35_Y_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_b_Y = pippenger_1_dataRam_1_1_io_rData_1_regNext_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_b_Y = pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_b_Y = pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_b_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_b_Z = stage1_inputData_1_delay_35_Z_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_b_Z = pippenger_1_dataRam_1_1_io_rData_1_regNext_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_b_Z = pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_b_Z = pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_b_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_b_T = stage1_inputData_1_delay_35_T_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_b_T = pippenger_1_dataRam_1_1_io_rData_1_regNext_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_b_T = pippenger_1_dataRam_1_1_io_rData_1_regNext_T_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_b_T = pippenger_1_dataRam_1_1_io_rData_1_regNext_T_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_1_io_dataIn_1_payload_address = 16'bxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_1_io_dataIn_1_payload_address = stage1_inputAddress_1_delay_35;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_1_io_dataIn_1_payload_address = _zz_io_dataIn_1_payload_address_59;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_1_io_dataIn_1_payload_address = {_zz_io_dataIn_1_payload_address_119,12'h001};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        fifo_1_io_dataIn_1_payload_address = 16'h0001;
      end
      default : begin
      end
    endcase
  end

  assign io_dataOut_valid = outputValid;
  assign io_dataOut_payload_X = pAddPort_0_s_regNext_X;
  assign io_dataOut_payload_Y = pAddPort_0_s_regNext_Y;
  assign io_dataOut_payload_Z = pAddPort_0_s_regNext_Z;
  assign io_dataOut_payload_T = pAddPort_0_s_regNext_T;
  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    flushing_flushCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
        flushing_flushCnt_willIncrement = 1'b1;
      end
    endcase
  end

  assign flushing_flushCnt_willClear = 1'b0;
  assign flushing_flushCnt_willOverflow = (flushing_flushCnt_willOverflowIfInc && flushing_flushCnt_willIncrement);
  always @(*) begin
    if(flushing_flushCnt_willOverflow) begin
      flushing_flushCnt_valueNext = 16'h0;
    end else begin
      flushing_flushCnt_valueNext = (flushing_flushCnt_value + _zz_flushing_flushCnt_valueNext);
    end
    if(flushing_flushCnt_willClear) begin
      flushing_flushCnt_valueNext = 16'h0;
    end
  end

  always @(*) begin
    stage1_NCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          if(dataInBuffer_bufferOut_valid) begin
            if(stage1_GCnt_willOverflowIfInc) begin
              stage1_NCnt_willIncrement = 1'b1;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stage1_NCnt_willClear = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          if(dataInBuffer_bufferOut_valid) begin
            if(stage1_GCnt_willOverflowIfInc) begin
              if(dataInBuffer_bufferOut_payload_last) begin
                stage1_NCnt_willClear = 1'b1;
              end
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage1_NCnt_willOverflow = (stage1_NCnt_willOverflowIfInc && stage1_NCnt_willIncrement);
  always @(*) begin
    stage1_NCnt_valueNext = (stage1_NCnt_value + _zz_stage1_NCnt_valueNext);
    if(stage1_NCnt_willClear) begin
      stage1_NCnt_valueNext = 32'h0;
    end
  end

  always @(*) begin
    stage1_GCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          if(dataInBuffer_bufferOut_valid) begin
            stage1_GCnt_willIncrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage1_GCnt_willClear = 1'b0;
  assign stage1_GCnt_willOverflow = (stage1_GCnt_willOverflowIfInc && stage1_GCnt_willIncrement);
  always @(*) begin
    if(stage1_GCnt_willOverflow) begin
      stage1_GCnt_valueNext = 4'b0000;
    end else begin
      stage1_GCnt_valueNext = (stage1_GCnt_value + _zz_stage1_GCnt_valueNext);
    end
    if(stage1_GCnt_willClear) begin
      stage1_GCnt_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    stage1_emptyCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(!when_Pippenger_l153) begin
          if(!when_Pippenger_l168) begin
            stage1_emptyCnt_willIncrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stage1_emptyCnt_willClear = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(!when_Pippenger_l153) begin
          if(when_Pippenger_l168) begin
            stage1_emptyCnt_willClear = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage1_emptyCnt_willOverflow = (stage1_emptyCnt_willOverflowIfInc && stage1_emptyCnt_willIncrement);
  always @(*) begin
    if(stage1_emptyCnt_willOverflow) begin
      stage1_emptyCnt_valueNext = 9'h0;
    end else begin
      stage1_emptyCnt_valueNext = (stage1_emptyCnt_value + _zz_stage1_emptyCnt_valueNext);
    end
    if(stage1_emptyCnt_willClear) begin
      stage1_emptyCnt_valueNext = 9'h0;
    end
  end

  assign _zz_stage1_inputBarrelID_0 = dataInBuffer_bufferOut_payload_fragment_K[25:0];
  assign stage1_inputBarrelID_0 = ({1'b0,_zz_stage1_inputBarrelID_0[12 : 0]} + _zz_stage1_inputBarrelID_0_1);
  assign stage1_inputBarrelID_1 = ({1'b0,_zz_stage1_inputBarrelID_0[25 : 13]} + _zz_stage1_inputBarrelID_1);
  assign _zz_stage1_inputBarrelIDAbs_0 = _zz__zz_stage1_inputBarrelIDAbs_0;
  assign stage1_inputBarrelIDAbs_0 = _zz_stage1_inputBarrelIDAbs_0_1[11:0];
  assign _zz_stage1_inputBarrelIDAbs_1 = _zz__zz_stage1_inputBarrelIDAbs_1;
  assign stage1_inputBarrelIDAbs_1 = _zz_stage1_inputBarrelIDAbs_1_1[11:0];
  assign stage1_inputData_0_X = (_zz_stage1_inputData_0_X_5 ? pNegPort_n_X : dataInBuffer_bufferOut_payload_fragment_P_delay_6_X);
  assign stage1_inputData_0_Y = (_zz_stage1_inputData_0_X_5 ? pNegPort_n_Y : dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y);
  assign stage1_inputData_0_Z = (_zz_stage1_inputData_0_X_5 ? pNegPort_n_Z : dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z);
  assign stage1_inputData_0_T = (_zz_stage1_inputData_0_X_5 ? pNegPort_n_T : dataInBuffer_bufferOut_payload_fragment_P_delay_6_T);
  assign stage1_inputData_1_X = (_zz_stage1_inputData_1_X_5 ? pNegPort_n_X : dataInBuffer_bufferOut_payload_fragment_P_delay_6_X_1);
  assign stage1_inputData_1_Y = (_zz_stage1_inputData_1_X_5 ? pNegPort_n_Y : dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y_1);
  assign stage1_inputData_1_Z = (_zz_stage1_inputData_1_X_5 ? pNegPort_n_Z : dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z_1);
  assign stage1_inputData_1_T = (_zz_stage1_inputData_1_X_5 ? pNegPort_n_T : dataInBuffer_bufferOut_payload_fragment_P_delay_6_T_1);
  assign pAddPort_0_a_X = fifo_0_io_dataOut_payload_a_X;
  assign pAddPort_0_a_Y = fifo_0_io_dataOut_payload_a_Y;
  assign pAddPort_0_a_Z = fifo_0_io_dataOut_payload_a_Z;
  assign pAddPort_0_a_T = fifo_0_io_dataOut_payload_a_T;
  assign pAddPort_1_a_X = fifo_1_io_dataOut_payload_a_X;
  assign pAddPort_1_a_Y = fifo_1_io_dataOut_payload_a_Y;
  assign pAddPort_1_a_Z = fifo_1_io_dataOut_payload_a_Z;
  assign pAddPort_1_a_T = fifo_1_io_dataOut_payload_a_T;
  assign pAddPort_0_b_X = fifo_0_io_dataOut_payload_b_X;
  assign pAddPort_0_b_Y = fifo_0_io_dataOut_payload_b_Y;
  assign pAddPort_0_b_Z = fifo_0_io_dataOut_payload_b_Z;
  assign pAddPort_0_b_T = fifo_0_io_dataOut_payload_b_T;
  assign pAddPort_1_b_X = fifo_1_io_dataOut_payload_b_X;
  assign pAddPort_1_b_Y = fifo_1_io_dataOut_payload_b_Y;
  assign pAddPort_1_b_Z = fifo_1_io_dataOut_payload_b_Z;
  assign pAddPort_1_b_T = fifo_1_io_dataOut_payload_b_T;
  assign pNegPort_a_X = dataInBuffer_bufferOut_payload_fragment_P_X;
  assign pNegPort_a_Y = dataInBuffer_bufferOut_payload_fragment_P_Y;
  assign pNegPort_a_Z = dataInBuffer_bufferOut_payload_fragment_P_Z;
  assign pNegPort_a_T = dataInBuffer_bufferOut_payload_fragment_P_T;
  assign shiftRegs_validIn_0 = fifo_0_io_dataOut_valid;
  assign shiftRegs_validIn_1 = fifo_1_io_dataOut_valid;
  assign shiftRegs_addressIn_0 = fifo_0_io_dataOut_payload_address;
  assign shiftRegs_addressIn_1 = fifo_1_io_dataOut_payload_address;
  always @(*) begin
    stage2_wCnt_willDecrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(!when_Pippenger_l207) begin
          if(stage2_waitCnt_willOverflowIfInc) begin
            stage2_wCnt_willDecrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage2_wCnt_willClear = 1'b0;
  assign stage2_wCnt_willUnderflow = (stage2_wCnt_willUnderflowIfDec && stage2_wCnt_willDecrement);
  always @(*) begin
    stage2_wCnt_valueNext = (stage2_wCnt_value - _zz_stage2_wCnt_valueNext);
    if(stage2_wCnt_willClear) begin
      stage2_wCnt_valueNext = 12'hfff;
    end
  end

  always @(*) begin
    stage2_GCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(when_Pippenger_l207) begin
          if(stage2_calCnt_willUnderflowIfDec) begin
            stage2_GCnt_willIncrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage2_GCnt_willClear = 1'b0;
  assign stage2_GCnt_willOverflow = (stage2_GCnt_willOverflowIfInc && stage2_GCnt_willIncrement);
  always @(*) begin
    if(stage2_GCnt_willOverflow) begin
      stage2_GCnt_valueNext = 4'b0000;
    end else begin
      stage2_GCnt_valueNext = (stage2_GCnt_value + _zz_stage2_GCnt_valueNext);
    end
    if(stage2_GCnt_willClear) begin
      stage2_GCnt_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    stage2_calCnt_willDecrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(when_Pippenger_l207) begin
          stage2_calCnt_willDecrement = 1'b1;
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage2_calCnt_willClear = 1'b0;
  assign stage2_calCnt_willUnderflow = (stage2_calCnt_willUnderflowIfDec && stage2_calCnt_willDecrement);
  always @(*) begin
    if(stage2_calCnt_willUnderflow) begin
      stage2_calCnt_valueNext = 2'b10;
    end else begin
      stage2_calCnt_valueNext = (stage2_calCnt_value - _zz_stage2_calCnt_valueNext);
    end
    if(stage2_calCnt_willClear) begin
      stage2_calCnt_valueNext = 2'b10;
    end
  end

  always @(*) begin
    stage2_waitCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(!when_Pippenger_l207) begin
          stage2_waitCnt_willIncrement = 1'b1;
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage2_waitCnt_willClear = 1'b0;
  assign stage2_waitCnt_willOverflow = (stage2_waitCnt_willOverflowIfInc && stage2_waitCnt_willIncrement);
  always @(*) begin
    if(stage2_waitCnt_willOverflow) begin
      stage2_waitCnt_valueNext = 9'h0;
    end else begin
      stage2_waitCnt_valueNext = (stage2_waitCnt_value + _zz_stage2_waitCnt_valueNext);
    end
    if(stage2_waitCnt_willClear) begin
      stage2_waitCnt_valueNext = 9'h0;
    end
  end

  always @(*) begin
    stage3_GCnt_willDecrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(!when_Pippenger_l249) begin
          if(stage3_addWaitCnt_willOverflowIfInc) begin
            stage3_GCnt_willDecrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage3_GCnt_willClear = 1'b0;
  assign stage3_GCnt_willUnderflow = (stage3_GCnt_willUnderflowIfDec && stage3_GCnt_willDecrement);
  always @(*) begin
    if(stage3_GCnt_willUnderflow) begin
      stage3_GCnt_valueNext = 4'b1001;
    end else begin
      stage3_GCnt_valueNext = (stage3_GCnt_value - _zz_stage3_GCnt_valueNext);
    end
    if(stage3_GCnt_willClear) begin
      stage3_GCnt_valueNext = 4'b1001;
    end
  end

  always @(*) begin
    stage3_doubleCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(when_Pippenger_l249) begin
          if(stage3_doubleWaitCnt_willOverflowIfInc) begin
            stage3_doubleCnt_willIncrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage3_doubleCnt_willClear = 1'b0;
  assign stage3_doubleCnt_willOverflow = (stage3_doubleCnt_willOverflowIfInc && stage3_doubleCnt_willIncrement);
  always @(*) begin
    if(stage3_doubleCnt_willOverflow) begin
      stage3_doubleCnt_valueNext = 5'h0;
    end else begin
      stage3_doubleCnt_valueNext = (stage3_doubleCnt_value + _zz_stage3_doubleCnt_valueNext);
    end
    if(stage3_doubleCnt_willClear) begin
      stage3_doubleCnt_valueNext = 5'h0;
    end
  end

  always @(*) begin
    stage3_doubleWaitCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(when_Pippenger_l249) begin
          stage3_doubleWaitCnt_willIncrement = 1'b1;
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage3_doubleWaitCnt_willClear = 1'b0;
  assign stage3_doubleWaitCnt_willOverflow = (stage3_doubleWaitCnt_willOverflowIfInc && stage3_doubleWaitCnt_willIncrement);
  always @(*) begin
    if(stage3_doubleWaitCnt_willOverflow) begin
      stage3_doubleWaitCnt_valueNext = 9'h0;
    end else begin
      stage3_doubleWaitCnt_valueNext = (stage3_doubleWaitCnt_value + _zz_stage3_doubleWaitCnt_valueNext);
    end
    if(stage3_doubleWaitCnt_willClear) begin
      stage3_doubleWaitCnt_valueNext = 9'h0;
    end
  end

  always @(*) begin
    stage3_addWaitCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(!when_Pippenger_l249) begin
          stage3_addWaitCnt_willIncrement = 1'b1;
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage3_addWaitCnt_willClear = 1'b0;
  assign stage3_addWaitCnt_willOverflow = (stage3_addWaitCnt_willOverflowIfInc && stage3_addWaitCnt_willIncrement);
  always @(*) begin
    if(stage3_addWaitCnt_willOverflow) begin
      stage3_addWaitCnt_valueNext = 9'h0;
    end else begin
      stage3_addWaitCnt_valueNext = (stage3_addWaitCnt_value + _zz_stage3_addWaitCnt_valueNext);
    end
    if(stage3_addWaitCnt_willClear) begin
      stage3_addWaitCnt_valueNext = 9'h0;
    end
  end

  always @(*) begin
    stage3Final_doubleCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        if(when_Pippenger_l306) begin
          if(stage3Final_doubleWaitCnt_willOverflowIfInc) begin
            stage3Final_doubleCnt_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign stage3Final_doubleCnt_willClear = 1'b0;
  assign stage3Final_doubleCnt_willOverflow = (stage3Final_doubleCnt_willOverflowIfInc && stage3Final_doubleCnt_willIncrement);
  always @(*) begin
    if(stage3Final_doubleCnt_willOverflow) begin
      stage3Final_doubleCnt_valueNext = 4'b0000;
    end else begin
      stage3Final_doubleCnt_valueNext = (stage3Final_doubleCnt_value + _zz_stage3Final_doubleCnt_valueNext);
    end
    if(stage3Final_doubleCnt_willClear) begin
      stage3Final_doubleCnt_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    stage3Final_doubleWaitCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        if(when_Pippenger_l306) begin
          stage3Final_doubleWaitCnt_willIncrement = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign stage3Final_doubleWaitCnt_willClear = 1'b0;
  assign stage3Final_doubleWaitCnt_willOverflow = (stage3Final_doubleWaitCnt_willOverflowIfInc && stage3Final_doubleWaitCnt_willIncrement);
  always @(*) begin
    if(stage3Final_doubleWaitCnt_willOverflow) begin
      stage3Final_doubleWaitCnt_valueNext = 9'h0;
    end else begin
      stage3Final_doubleWaitCnt_valueNext = (stage3Final_doubleWaitCnt_value + _zz_stage3Final_doubleWaitCnt_valueNext);
    end
    if(stage3Final_doubleWaitCnt_willClear) begin
      stage3Final_doubleWaitCnt_valueNext = 9'h0;
    end
  end

  always @(*) begin
    stage3Final_addWaitCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        if(!when_Pippenger_l306) begin
          stage3Final_addWaitCnt_willIncrement = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign stage3Final_addWaitCnt_willClear = 1'b0;
  assign stage3Final_addWaitCnt_willOverflow = (stage3Final_addWaitCnt_willOverflowIfInc && stage3Final_addWaitCnt_willIncrement);
  always @(*) begin
    if(stage3Final_addWaitCnt_willOverflow) begin
      stage3Final_addWaitCnt_valueNext = 9'h0;
    end else begin
      stage3Final_addWaitCnt_valueNext = (stage3Final_addWaitCnt_value + _zz_stage3Final_addWaitCnt_valueNext);
    end
    if(stage3Final_addWaitCnt_willClear) begin
      stage3Final_addWaitCnt_valueNext = 9'h0;
    end
  end

  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(!when_Pippenger_l153) begin
          if(!when_Pippenger_l168) begin
            if(stage1_emptyCnt_willOverflowIfInc) begin
              fsm_stateNext = fsm_enumDef_stage2;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(!when_Pippenger_l207) begin
          if(stage2_waitCnt_willOverflowIfInc) begin
            if(stage2_wCnt_willUnderflowIfDec) begin
              fsm_stateNext = fsm_enumDef_stage3;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(!when_Pippenger_l249) begin
          if(stage3_addWaitCnt_willOverflowIfInc) begin
            if(stage3_GCnt_willUnderflowIfDec) begin
              fsm_stateNext = fsm_enumDef_stage3Final;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
        if(!when_Pippenger_l306) begin
          if(stage3Final_addWaitCnt_willOverflowIfInc) begin
            if(when_Pippenger_l319) begin
              fsm_stateNext = fsm_enumDef_stage1;
            end
          end
        end
      end
      default : begin
        if(flushing_flushCnt_willOverflowIfInc) begin
          fsm_stateNext = fsm_enumDef_stage1;
        end
      end
    endcase
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_flushing;
    end
  end

  assign when_Pippenger_l153 = (! stage1_waitReg);
  assign when_Pippenger_l168 = ({fifo_1_io_dataOut_valid,fifo_0_io_dataOut_valid} != 2'b00);
  assign when_Pippenger_l207 = (! stage2_waitReg);
  assign when_Pippenger_l249 = (! stage3_addReg);
  assign when_Pippenger_l306 = (! stage3Final_addReg);
  assign when_Pippenger_l319 = stage3Final_pAddShr[0];
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      dataInBuffer_validReg <= 1'b0;
      shiftRegs_validIn_delay_1_0 <= 1'b0;
      shiftRegs_validIn_delay_1_1 <= 1'b0;
      shiftRegs_validIn_delay_2_0 <= 1'b0;
      shiftRegs_validIn_delay_2_1 <= 1'b0;
      shiftRegs_validIn_delay_3_0 <= 1'b0;
      shiftRegs_validIn_delay_3_1 <= 1'b0;
      shiftRegs_validIn_delay_4_0 <= 1'b0;
      shiftRegs_validIn_delay_4_1 <= 1'b0;
      shiftRegs_validIn_delay_5_0 <= 1'b0;
      shiftRegs_validIn_delay_5_1 <= 1'b0;
      shiftRegs_validIn_delay_6_0 <= 1'b0;
      shiftRegs_validIn_delay_6_1 <= 1'b0;
      shiftRegs_validIn_delay_7_0 <= 1'b0;
      shiftRegs_validIn_delay_7_1 <= 1'b0;
      shiftRegs_validIn_delay_8_0 <= 1'b0;
      shiftRegs_validIn_delay_8_1 <= 1'b0;
      shiftRegs_validIn_delay_9_0 <= 1'b0;
      shiftRegs_validIn_delay_9_1 <= 1'b0;
      shiftRegs_validIn_delay_10_0 <= 1'b0;
      shiftRegs_validIn_delay_10_1 <= 1'b0;
      shiftRegs_validIn_delay_11_0 <= 1'b0;
      shiftRegs_validIn_delay_11_1 <= 1'b0;
      shiftRegs_validIn_delay_12_0 <= 1'b0;
      shiftRegs_validIn_delay_12_1 <= 1'b0;
      shiftRegs_validIn_delay_13_0 <= 1'b0;
      shiftRegs_validIn_delay_13_1 <= 1'b0;
      shiftRegs_validIn_delay_14_0 <= 1'b0;
      shiftRegs_validIn_delay_14_1 <= 1'b0;
      shiftRegs_validIn_delay_15_0 <= 1'b0;
      shiftRegs_validIn_delay_15_1 <= 1'b0;
      shiftRegs_validIn_delay_16_0 <= 1'b0;
      shiftRegs_validIn_delay_16_1 <= 1'b0;
      shiftRegs_validIn_delay_17_0 <= 1'b0;
      shiftRegs_validIn_delay_17_1 <= 1'b0;
      shiftRegs_validIn_delay_18_0 <= 1'b0;
      shiftRegs_validIn_delay_18_1 <= 1'b0;
      shiftRegs_validIn_delay_19_0 <= 1'b0;
      shiftRegs_validIn_delay_19_1 <= 1'b0;
      shiftRegs_validIn_delay_20_0 <= 1'b0;
      shiftRegs_validIn_delay_20_1 <= 1'b0;
      shiftRegs_validIn_delay_21_0 <= 1'b0;
      shiftRegs_validIn_delay_21_1 <= 1'b0;
      shiftRegs_validIn_delay_22_0 <= 1'b0;
      shiftRegs_validIn_delay_22_1 <= 1'b0;
      shiftRegs_validIn_delay_23_0 <= 1'b0;
      shiftRegs_validIn_delay_23_1 <= 1'b0;
      shiftRegs_validIn_delay_24_0 <= 1'b0;
      shiftRegs_validIn_delay_24_1 <= 1'b0;
      shiftRegs_validIn_delay_25_0 <= 1'b0;
      shiftRegs_validIn_delay_25_1 <= 1'b0;
      shiftRegs_validIn_delay_26_0 <= 1'b0;
      shiftRegs_validIn_delay_26_1 <= 1'b0;
      shiftRegs_validIn_delay_27_0 <= 1'b0;
      shiftRegs_validIn_delay_27_1 <= 1'b0;
      shiftRegs_validIn_delay_28_0 <= 1'b0;
      shiftRegs_validIn_delay_28_1 <= 1'b0;
      shiftRegs_validIn_delay_29_0 <= 1'b0;
      shiftRegs_validIn_delay_29_1 <= 1'b0;
      shiftRegs_validIn_delay_30_0 <= 1'b0;
      shiftRegs_validIn_delay_30_1 <= 1'b0;
      shiftRegs_validIn_delay_31_0 <= 1'b0;
      shiftRegs_validIn_delay_31_1 <= 1'b0;
      shiftRegs_validIn_delay_32_0 <= 1'b0;
      shiftRegs_validIn_delay_32_1 <= 1'b0;
      shiftRegs_validIn_delay_33_0 <= 1'b0;
      shiftRegs_validIn_delay_33_1 <= 1'b0;
      shiftRegs_validIn_delay_34_0 <= 1'b0;
      shiftRegs_validIn_delay_34_1 <= 1'b0;
      shiftRegs_validIn_delay_35_0 <= 1'b0;
      shiftRegs_validIn_delay_35_1 <= 1'b0;
      shiftRegs_validIn_delay_36_0 <= 1'b0;
      shiftRegs_validIn_delay_36_1 <= 1'b0;
      shiftRegs_validIn_delay_37_0 <= 1'b0;
      shiftRegs_validIn_delay_37_1 <= 1'b0;
      shiftRegs_validIn_delay_38_0 <= 1'b0;
      shiftRegs_validIn_delay_38_1 <= 1'b0;
      shiftRegs_validIn_delay_39_0 <= 1'b0;
      shiftRegs_validIn_delay_39_1 <= 1'b0;
      shiftRegs_validIn_delay_40_0 <= 1'b0;
      shiftRegs_validIn_delay_40_1 <= 1'b0;
      shiftRegs_validIn_delay_41_0 <= 1'b0;
      shiftRegs_validIn_delay_41_1 <= 1'b0;
      shiftRegs_validIn_delay_42_0 <= 1'b0;
      shiftRegs_validIn_delay_42_1 <= 1'b0;
      shiftRegs_validIn_delay_43_0 <= 1'b0;
      shiftRegs_validIn_delay_43_1 <= 1'b0;
      shiftRegs_validIn_delay_44_0 <= 1'b0;
      shiftRegs_validIn_delay_44_1 <= 1'b0;
      shiftRegs_validIn_delay_45_0 <= 1'b0;
      shiftRegs_validIn_delay_45_1 <= 1'b0;
      shiftRegs_validIn_delay_46_0 <= 1'b0;
      shiftRegs_validIn_delay_46_1 <= 1'b0;
      shiftRegs_validIn_delay_47_0 <= 1'b0;
      shiftRegs_validIn_delay_47_1 <= 1'b0;
      shiftRegs_validIn_delay_48_0 <= 1'b0;
      shiftRegs_validIn_delay_48_1 <= 1'b0;
      shiftRegs_validIn_delay_49_0 <= 1'b0;
      shiftRegs_validIn_delay_49_1 <= 1'b0;
      shiftRegs_validIn_delay_50_0 <= 1'b0;
      shiftRegs_validIn_delay_50_1 <= 1'b0;
      shiftRegs_validIn_delay_51_0 <= 1'b0;
      shiftRegs_validIn_delay_51_1 <= 1'b0;
      shiftRegs_validIn_delay_52_0 <= 1'b0;
      shiftRegs_validIn_delay_52_1 <= 1'b0;
      shiftRegs_validIn_delay_53_0 <= 1'b0;
      shiftRegs_validIn_delay_53_1 <= 1'b0;
      shiftRegs_validIn_delay_54_0 <= 1'b0;
      shiftRegs_validIn_delay_54_1 <= 1'b0;
      shiftRegs_validIn_delay_55_0 <= 1'b0;
      shiftRegs_validIn_delay_55_1 <= 1'b0;
      shiftRegs_validIn_delay_56_0 <= 1'b0;
      shiftRegs_validIn_delay_56_1 <= 1'b0;
      shiftRegs_validIn_delay_57_0 <= 1'b0;
      shiftRegs_validIn_delay_57_1 <= 1'b0;
      shiftRegs_validIn_delay_58_0 <= 1'b0;
      shiftRegs_validIn_delay_58_1 <= 1'b0;
      shiftRegs_validIn_delay_59_0 <= 1'b0;
      shiftRegs_validIn_delay_59_1 <= 1'b0;
      shiftRegs_validIn_delay_60_0 <= 1'b0;
      shiftRegs_validIn_delay_60_1 <= 1'b0;
      shiftRegs_validIn_delay_61_0 <= 1'b0;
      shiftRegs_validIn_delay_61_1 <= 1'b0;
      shiftRegs_validIn_delay_62_0 <= 1'b0;
      shiftRegs_validIn_delay_62_1 <= 1'b0;
      shiftRegs_validIn_delay_63_0 <= 1'b0;
      shiftRegs_validIn_delay_63_1 <= 1'b0;
      shiftRegs_validIn_delay_64_0 <= 1'b0;
      shiftRegs_validIn_delay_64_1 <= 1'b0;
      shiftRegs_validIn_delay_65_0 <= 1'b0;
      shiftRegs_validIn_delay_65_1 <= 1'b0;
      shiftRegs_validIn_delay_66_0 <= 1'b0;
      shiftRegs_validIn_delay_66_1 <= 1'b0;
      shiftRegs_validIn_delay_67_0 <= 1'b0;
      shiftRegs_validIn_delay_67_1 <= 1'b0;
      shiftRegs_validIn_delay_68_0 <= 1'b0;
      shiftRegs_validIn_delay_68_1 <= 1'b0;
      shiftRegs_validIn_delay_69_0 <= 1'b0;
      shiftRegs_validIn_delay_69_1 <= 1'b0;
      shiftRegs_validIn_delay_70_0 <= 1'b0;
      shiftRegs_validIn_delay_70_1 <= 1'b0;
      shiftRegs_validIn_delay_71_0 <= 1'b0;
      shiftRegs_validIn_delay_71_1 <= 1'b0;
      shiftRegs_validIn_delay_72_0 <= 1'b0;
      shiftRegs_validIn_delay_72_1 <= 1'b0;
      shiftRegs_validIn_delay_73_0 <= 1'b0;
      shiftRegs_validIn_delay_73_1 <= 1'b0;
      shiftRegs_validIn_delay_74_0 <= 1'b0;
      shiftRegs_validIn_delay_74_1 <= 1'b0;
      shiftRegs_validIn_delay_75_0 <= 1'b0;
      shiftRegs_validIn_delay_75_1 <= 1'b0;
      shiftRegs_validIn_delay_76_0 <= 1'b0;
      shiftRegs_validIn_delay_76_1 <= 1'b0;
      shiftRegs_validIn_delay_77_0 <= 1'b0;
      shiftRegs_validIn_delay_77_1 <= 1'b0;
      shiftRegs_validIn_delay_78_0 <= 1'b0;
      shiftRegs_validIn_delay_78_1 <= 1'b0;
      shiftRegs_validIn_delay_79_0 <= 1'b0;
      shiftRegs_validIn_delay_79_1 <= 1'b0;
      shiftRegs_validIn_delay_80_0 <= 1'b0;
      shiftRegs_validIn_delay_80_1 <= 1'b0;
      shiftRegs_validIn_delay_81_0 <= 1'b0;
      shiftRegs_validIn_delay_81_1 <= 1'b0;
      shiftRegs_validIn_delay_82_0 <= 1'b0;
      shiftRegs_validIn_delay_82_1 <= 1'b0;
      shiftRegs_validIn_delay_83_0 <= 1'b0;
      shiftRegs_validIn_delay_83_1 <= 1'b0;
      shiftRegs_validIn_delay_84_0 <= 1'b0;
      shiftRegs_validIn_delay_84_1 <= 1'b0;
      shiftRegs_validIn_delay_85_0 <= 1'b0;
      shiftRegs_validIn_delay_85_1 <= 1'b0;
      shiftRegs_validIn_delay_86_0 <= 1'b0;
      shiftRegs_validIn_delay_86_1 <= 1'b0;
      shiftRegs_validIn_delay_87_0 <= 1'b0;
      shiftRegs_validIn_delay_87_1 <= 1'b0;
      shiftRegs_validIn_delay_88_0 <= 1'b0;
      shiftRegs_validIn_delay_88_1 <= 1'b0;
      shiftRegs_validIn_delay_89_0 <= 1'b0;
      shiftRegs_validIn_delay_89_1 <= 1'b0;
      shiftRegs_validIn_delay_90_0 <= 1'b0;
      shiftRegs_validIn_delay_90_1 <= 1'b0;
      shiftRegs_validIn_delay_91_0 <= 1'b0;
      shiftRegs_validIn_delay_91_1 <= 1'b0;
      shiftRegs_validIn_delay_92_0 <= 1'b0;
      shiftRegs_validIn_delay_92_1 <= 1'b0;
      shiftRegs_validIn_delay_93_0 <= 1'b0;
      shiftRegs_validIn_delay_93_1 <= 1'b0;
      shiftRegs_validIn_delay_94_0 <= 1'b0;
      shiftRegs_validIn_delay_94_1 <= 1'b0;
      shiftRegs_validIn_delay_95_0 <= 1'b0;
      shiftRegs_validIn_delay_95_1 <= 1'b0;
      shiftRegs_validIn_delay_96_0 <= 1'b0;
      shiftRegs_validIn_delay_96_1 <= 1'b0;
      shiftRegs_validIn_delay_97_0 <= 1'b0;
      shiftRegs_validIn_delay_97_1 <= 1'b0;
      shiftRegs_validIn_delay_98_0 <= 1'b0;
      shiftRegs_validIn_delay_98_1 <= 1'b0;
      shiftRegs_validIn_delay_99_0 <= 1'b0;
      shiftRegs_validIn_delay_99_1 <= 1'b0;
      shiftRegs_validIn_delay_100_0 <= 1'b0;
      shiftRegs_validIn_delay_100_1 <= 1'b0;
      shiftRegs_validIn_delay_101_0 <= 1'b0;
      shiftRegs_validIn_delay_101_1 <= 1'b0;
      shiftRegs_validIn_delay_102_0 <= 1'b0;
      shiftRegs_validIn_delay_102_1 <= 1'b0;
      shiftRegs_validIn_delay_103_0 <= 1'b0;
      shiftRegs_validIn_delay_103_1 <= 1'b0;
      shiftRegs_validIn_delay_104_0 <= 1'b0;
      shiftRegs_validIn_delay_104_1 <= 1'b0;
      shiftRegs_validIn_delay_105_0 <= 1'b0;
      shiftRegs_validIn_delay_105_1 <= 1'b0;
      shiftRegs_validIn_delay_106_0 <= 1'b0;
      shiftRegs_validIn_delay_106_1 <= 1'b0;
      shiftRegs_validIn_delay_107_0 <= 1'b0;
      shiftRegs_validIn_delay_107_1 <= 1'b0;
      shiftRegs_validIn_delay_108_0 <= 1'b0;
      shiftRegs_validIn_delay_108_1 <= 1'b0;
      shiftRegs_validIn_delay_109_0 <= 1'b0;
      shiftRegs_validIn_delay_109_1 <= 1'b0;
      shiftRegs_validIn_delay_110_0 <= 1'b0;
      shiftRegs_validIn_delay_110_1 <= 1'b0;
      shiftRegs_validIn_delay_111_0 <= 1'b0;
      shiftRegs_validIn_delay_111_1 <= 1'b0;
      shiftRegs_validIn_delay_112_0 <= 1'b0;
      shiftRegs_validIn_delay_112_1 <= 1'b0;
      shiftRegs_validIn_delay_113_0 <= 1'b0;
      shiftRegs_validIn_delay_113_1 <= 1'b0;
      shiftRegs_validIn_delay_114_0 <= 1'b0;
      shiftRegs_validIn_delay_114_1 <= 1'b0;
      shiftRegs_validIn_delay_115_0 <= 1'b0;
      shiftRegs_validIn_delay_115_1 <= 1'b0;
      shiftRegs_validIn_delay_116_0 <= 1'b0;
      shiftRegs_validIn_delay_116_1 <= 1'b0;
      shiftRegs_validIn_delay_117_0 <= 1'b0;
      shiftRegs_validIn_delay_117_1 <= 1'b0;
      shiftRegs_validIn_delay_118_0 <= 1'b0;
      shiftRegs_validIn_delay_118_1 <= 1'b0;
      shiftRegs_validIn_delay_119_0 <= 1'b0;
      shiftRegs_validIn_delay_119_1 <= 1'b0;
      shiftRegs_validIn_delay_120_0 <= 1'b0;
      shiftRegs_validIn_delay_120_1 <= 1'b0;
      shiftRegs_validIn_delay_121_0 <= 1'b0;
      shiftRegs_validIn_delay_121_1 <= 1'b0;
      shiftRegs_validIn_delay_122_0 <= 1'b0;
      shiftRegs_validIn_delay_122_1 <= 1'b0;
      shiftRegs_validIn_delay_123_0 <= 1'b0;
      shiftRegs_validIn_delay_123_1 <= 1'b0;
      shiftRegs_validIn_delay_124_0 <= 1'b0;
      shiftRegs_validIn_delay_124_1 <= 1'b0;
      shiftRegs_validIn_delay_125_0 <= 1'b0;
      shiftRegs_validIn_delay_125_1 <= 1'b0;
      shiftRegs_validIn_delay_126_0 <= 1'b0;
      shiftRegs_validIn_delay_126_1 <= 1'b0;
      shiftRegs_validIn_delay_127_0 <= 1'b0;
      shiftRegs_validIn_delay_127_1 <= 1'b0;
      shiftRegs_validIn_delay_128_0 <= 1'b0;
      shiftRegs_validIn_delay_128_1 <= 1'b0;
      shiftRegs_validIn_delay_129_0 <= 1'b0;
      shiftRegs_validIn_delay_129_1 <= 1'b0;
      shiftRegs_validIn_delay_130_0 <= 1'b0;
      shiftRegs_validIn_delay_130_1 <= 1'b0;
      shiftRegs_validIn_delay_131_0 <= 1'b0;
      shiftRegs_validIn_delay_131_1 <= 1'b0;
      shiftRegs_validIn_delay_132_0 <= 1'b0;
      shiftRegs_validIn_delay_132_1 <= 1'b0;
      shiftRegs_validIn_delay_133_0 <= 1'b0;
      shiftRegs_validIn_delay_133_1 <= 1'b0;
      shiftRegs_validIn_delay_134_0 <= 1'b0;
      shiftRegs_validIn_delay_134_1 <= 1'b0;
      shiftRegs_validIn_delay_135_0 <= 1'b0;
      shiftRegs_validIn_delay_135_1 <= 1'b0;
      shiftRegs_validIn_delay_136_0 <= 1'b0;
      shiftRegs_validIn_delay_136_1 <= 1'b0;
      shiftRegs_validIn_delay_137_0 <= 1'b0;
      shiftRegs_validIn_delay_137_1 <= 1'b0;
      shiftRegs_validIn_delay_138_0 <= 1'b0;
      shiftRegs_validIn_delay_138_1 <= 1'b0;
      shiftRegs_validIn_delay_139_0 <= 1'b0;
      shiftRegs_validIn_delay_139_1 <= 1'b0;
      shiftRegs_validIn_delay_140_0 <= 1'b0;
      shiftRegs_validIn_delay_140_1 <= 1'b0;
      shiftRegs_validIn_delay_141_0 <= 1'b0;
      shiftRegs_validIn_delay_141_1 <= 1'b0;
      shiftRegs_validIn_delay_142_0 <= 1'b0;
      shiftRegs_validIn_delay_142_1 <= 1'b0;
      shiftRegs_validIn_delay_143_0 <= 1'b0;
      shiftRegs_validIn_delay_143_1 <= 1'b0;
      shiftRegs_validIn_delay_144_0 <= 1'b0;
      shiftRegs_validIn_delay_144_1 <= 1'b0;
      shiftRegs_validIn_delay_145_0 <= 1'b0;
      shiftRegs_validIn_delay_145_1 <= 1'b0;
      shiftRegs_validIn_delay_146_0 <= 1'b0;
      shiftRegs_validIn_delay_146_1 <= 1'b0;
      shiftRegs_validIn_delay_147_0 <= 1'b0;
      shiftRegs_validIn_delay_147_1 <= 1'b0;
      shiftRegs_validIn_delay_148_0 <= 1'b0;
      shiftRegs_validIn_delay_148_1 <= 1'b0;
      shiftRegs_validIn_delay_149_0 <= 1'b0;
      shiftRegs_validIn_delay_149_1 <= 1'b0;
      shiftRegs_validIn_delay_150_0 <= 1'b0;
      shiftRegs_validIn_delay_150_1 <= 1'b0;
      shiftRegs_validIn_delay_151_0 <= 1'b0;
      shiftRegs_validIn_delay_151_1 <= 1'b0;
      shiftRegs_validIn_delay_152_0 <= 1'b0;
      shiftRegs_validIn_delay_152_1 <= 1'b0;
      shiftRegs_validIn_delay_153_0 <= 1'b0;
      shiftRegs_validIn_delay_153_1 <= 1'b0;
      shiftRegs_validIn_delay_154_0 <= 1'b0;
      shiftRegs_validIn_delay_154_1 <= 1'b0;
      shiftRegs_validIn_delay_155_0 <= 1'b0;
      shiftRegs_validIn_delay_155_1 <= 1'b0;
      shiftRegs_validIn_delay_156_0 <= 1'b0;
      shiftRegs_validIn_delay_156_1 <= 1'b0;
      shiftRegs_validIn_delay_157_0 <= 1'b0;
      shiftRegs_validIn_delay_157_1 <= 1'b0;
      shiftRegs_validIn_delay_158_0 <= 1'b0;
      shiftRegs_validIn_delay_158_1 <= 1'b0;
      shiftRegs_validIn_delay_159_0 <= 1'b0;
      shiftRegs_validIn_delay_159_1 <= 1'b0;
      shiftRegs_validIn_delay_160_0 <= 1'b0;
      shiftRegs_validIn_delay_160_1 <= 1'b0;
      shiftRegs_validIn_delay_161_0 <= 1'b0;
      shiftRegs_validIn_delay_161_1 <= 1'b0;
      shiftRegs_validIn_delay_162_0 <= 1'b0;
      shiftRegs_validIn_delay_162_1 <= 1'b0;
      shiftRegs_validIn_delay_163_0 <= 1'b0;
      shiftRegs_validIn_delay_163_1 <= 1'b0;
      shiftRegs_validIn_delay_164_0 <= 1'b0;
      shiftRegs_validIn_delay_164_1 <= 1'b0;
      shiftRegs_validIn_delay_165_0 <= 1'b0;
      shiftRegs_validIn_delay_165_1 <= 1'b0;
      shiftRegs_validIn_delay_166_0 <= 1'b0;
      shiftRegs_validIn_delay_166_1 <= 1'b0;
      shiftRegs_validIn_delay_167_0 <= 1'b0;
      shiftRegs_validIn_delay_167_1 <= 1'b0;
      shiftRegs_validIn_delay_168_0 <= 1'b0;
      shiftRegs_validIn_delay_168_1 <= 1'b0;
      shiftRegs_validIn_delay_169_0 <= 1'b0;
      shiftRegs_validIn_delay_169_1 <= 1'b0;
      shiftRegs_validIn_delay_170_0 <= 1'b0;
      shiftRegs_validIn_delay_170_1 <= 1'b0;
      shiftRegs_validIn_delay_171_0 <= 1'b0;
      shiftRegs_validIn_delay_171_1 <= 1'b0;
      shiftRegs_validIn_delay_172_0 <= 1'b0;
      shiftRegs_validIn_delay_172_1 <= 1'b0;
      shiftRegs_validIn_delay_173_0 <= 1'b0;
      shiftRegs_validIn_delay_173_1 <= 1'b0;
      shiftRegs_validIn_delay_174_0 <= 1'b0;
      shiftRegs_validIn_delay_174_1 <= 1'b0;
      shiftRegs_validIn_delay_175_0 <= 1'b0;
      shiftRegs_validIn_delay_175_1 <= 1'b0;
      shiftRegs_validIn_delay_176_0 <= 1'b0;
      shiftRegs_validIn_delay_176_1 <= 1'b0;
      shiftRegs_validIn_delay_177_0 <= 1'b0;
      shiftRegs_validIn_delay_177_1 <= 1'b0;
      shiftRegs_validIn_delay_178_0 <= 1'b0;
      shiftRegs_validIn_delay_178_1 <= 1'b0;
      shiftRegs_validIn_delay_179_0 <= 1'b0;
      shiftRegs_validIn_delay_179_1 <= 1'b0;
      shiftRegs_validIn_delay_180_0 <= 1'b0;
      shiftRegs_validIn_delay_180_1 <= 1'b0;
      shiftRegs_validIn_delay_181_0 <= 1'b0;
      shiftRegs_validIn_delay_181_1 <= 1'b0;
      shiftRegs_validIn_delay_182_0 <= 1'b0;
      shiftRegs_validIn_delay_182_1 <= 1'b0;
      shiftRegs_validIn_delay_183_0 <= 1'b0;
      shiftRegs_validIn_delay_183_1 <= 1'b0;
      shiftRegs_validIn_delay_184_0 <= 1'b0;
      shiftRegs_validIn_delay_184_1 <= 1'b0;
      shiftRegs_validIn_delay_185_0 <= 1'b0;
      shiftRegs_validIn_delay_185_1 <= 1'b0;
      shiftRegs_validIn_delay_186_0 <= 1'b0;
      shiftRegs_validIn_delay_186_1 <= 1'b0;
      shiftRegs_validIn_delay_187_0 <= 1'b0;
      shiftRegs_validIn_delay_187_1 <= 1'b0;
      shiftRegs_validIn_delay_188_0 <= 1'b0;
      shiftRegs_validIn_delay_188_1 <= 1'b0;
      shiftRegs_validIn_delay_189_0 <= 1'b0;
      shiftRegs_validIn_delay_189_1 <= 1'b0;
      shiftRegs_validIn_delay_190_0 <= 1'b0;
      shiftRegs_validIn_delay_190_1 <= 1'b0;
      shiftRegs_validIn_delay_191_0 <= 1'b0;
      shiftRegs_validIn_delay_191_1 <= 1'b0;
      shiftRegs_validIn_delay_192_0 <= 1'b0;
      shiftRegs_validIn_delay_192_1 <= 1'b0;
      shiftRegs_validIn_delay_193_0 <= 1'b0;
      shiftRegs_validIn_delay_193_1 <= 1'b0;
      shiftRegs_validIn_delay_194_0 <= 1'b0;
      shiftRegs_validIn_delay_194_1 <= 1'b0;
      shiftRegs_validIn_delay_195_0 <= 1'b0;
      shiftRegs_validIn_delay_195_1 <= 1'b0;
      shiftRegs_validIn_delay_196_0 <= 1'b0;
      shiftRegs_validIn_delay_196_1 <= 1'b0;
      shiftRegs_validIn_delay_197_0 <= 1'b0;
      shiftRegs_validIn_delay_197_1 <= 1'b0;
      shiftRegs_validIn_delay_198_0 <= 1'b0;
      shiftRegs_validIn_delay_198_1 <= 1'b0;
      shiftRegs_validIn_delay_199_0 <= 1'b0;
      shiftRegs_validIn_delay_199_1 <= 1'b0;
      shiftRegs_validIn_delay_200_0 <= 1'b0;
      shiftRegs_validIn_delay_200_1 <= 1'b0;
      shiftRegs_validIn_delay_201_0 <= 1'b0;
      shiftRegs_validIn_delay_201_1 <= 1'b0;
      shiftRegs_validIn_delay_202_0 <= 1'b0;
      shiftRegs_validIn_delay_202_1 <= 1'b0;
      shiftRegs_validIn_delay_203_0 <= 1'b0;
      shiftRegs_validIn_delay_203_1 <= 1'b0;
      shiftRegs_validIn_delay_204_0 <= 1'b0;
      shiftRegs_validIn_delay_204_1 <= 1'b0;
      shiftRegs_validIn_delay_205_0 <= 1'b0;
      shiftRegs_validIn_delay_205_1 <= 1'b0;
      shiftRegs_validIn_delay_206_0 <= 1'b0;
      shiftRegs_validIn_delay_206_1 <= 1'b0;
      shiftRegs_validIn_delay_207_0 <= 1'b0;
      shiftRegs_validIn_delay_207_1 <= 1'b0;
      shiftRegs_validIn_delay_208_0 <= 1'b0;
      shiftRegs_validIn_delay_208_1 <= 1'b0;
      shiftRegs_validIn_delay_209_0 <= 1'b0;
      shiftRegs_validIn_delay_209_1 <= 1'b0;
      shiftRegs_validIn_delay_210_0 <= 1'b0;
      shiftRegs_validIn_delay_210_1 <= 1'b0;
      shiftRegs_validIn_delay_211_0 <= 1'b0;
      shiftRegs_validIn_delay_211_1 <= 1'b0;
      shiftRegs_validIn_delay_212_0 <= 1'b0;
      shiftRegs_validIn_delay_212_1 <= 1'b0;
      shiftRegs_validIn_delay_213_0 <= 1'b0;
      shiftRegs_validIn_delay_213_1 <= 1'b0;
      shiftRegs_validIn_delay_214_0 <= 1'b0;
      shiftRegs_validIn_delay_214_1 <= 1'b0;
      shiftRegs_validIn_delay_215_0 <= 1'b0;
      shiftRegs_validIn_delay_215_1 <= 1'b0;
      shiftRegs_validIn_delay_216_0 <= 1'b0;
      shiftRegs_validIn_delay_216_1 <= 1'b0;
      shiftRegs_validIn_delay_217_0 <= 1'b0;
      shiftRegs_validIn_delay_217_1 <= 1'b0;
      shiftRegs_validIn_delay_218_0 <= 1'b0;
      shiftRegs_validIn_delay_218_1 <= 1'b0;
      shiftRegs_validIn_delay_219_0 <= 1'b0;
      shiftRegs_validIn_delay_219_1 <= 1'b0;
      shiftRegs_validIn_delay_220_0 <= 1'b0;
      shiftRegs_validIn_delay_220_1 <= 1'b0;
      shiftRegs_validIn_delay_221_0 <= 1'b0;
      shiftRegs_validIn_delay_221_1 <= 1'b0;
      shiftRegs_validIn_delay_222_0 <= 1'b0;
      shiftRegs_validIn_delay_222_1 <= 1'b0;
      shiftRegs_validIn_delay_223_0 <= 1'b0;
      shiftRegs_validIn_delay_223_1 <= 1'b0;
      shiftRegs_validIn_delay_224_0 <= 1'b0;
      shiftRegs_validIn_delay_224_1 <= 1'b0;
      shiftRegs_validIn_delay_225_0 <= 1'b0;
      shiftRegs_validIn_delay_225_1 <= 1'b0;
      shiftRegs_validIn_delay_226_0 <= 1'b0;
      shiftRegs_validIn_delay_226_1 <= 1'b0;
      shiftRegs_validIn_delay_227_0 <= 1'b0;
      shiftRegs_validIn_delay_227_1 <= 1'b0;
      shiftRegs_validIn_delay_228_0 <= 1'b0;
      shiftRegs_validIn_delay_228_1 <= 1'b0;
      shiftRegs_validIn_delay_229_0 <= 1'b0;
      shiftRegs_validIn_delay_229_1 <= 1'b0;
      shiftRegs_validIn_delay_230_0 <= 1'b0;
      shiftRegs_validIn_delay_230_1 <= 1'b0;
      shiftRegs_validIn_delay_231_0 <= 1'b0;
      shiftRegs_validIn_delay_231_1 <= 1'b0;
      shiftRegs_validIn_delay_232_0 <= 1'b0;
      shiftRegs_validIn_delay_232_1 <= 1'b0;
      shiftRegs_validIn_delay_233_0 <= 1'b0;
      shiftRegs_validIn_delay_233_1 <= 1'b0;
      shiftRegs_validIn_delay_234_0 <= 1'b0;
      shiftRegs_validIn_delay_234_1 <= 1'b0;
      shiftRegs_validIn_delay_235_0 <= 1'b0;
      shiftRegs_validIn_delay_235_1 <= 1'b0;
      shiftRegs_validIn_delay_236_0 <= 1'b0;
      shiftRegs_validIn_delay_236_1 <= 1'b0;
      shiftRegs_validIn_delay_237_0 <= 1'b0;
      shiftRegs_validIn_delay_237_1 <= 1'b0;
      shiftRegs_validIn_delay_238_0 <= 1'b0;
      shiftRegs_validIn_delay_238_1 <= 1'b0;
      shiftRegs_validIn_delay_239_0 <= 1'b0;
      shiftRegs_validIn_delay_239_1 <= 1'b0;
      shiftRegs_validIn_delay_240_0 <= 1'b0;
      shiftRegs_validIn_delay_240_1 <= 1'b0;
      shiftRegs_validIn_delay_241_0 <= 1'b0;
      shiftRegs_validIn_delay_241_1 <= 1'b0;
      shiftRegs_validIn_delay_242_0 <= 1'b0;
      shiftRegs_validIn_delay_242_1 <= 1'b0;
      shiftRegs_validIn_delay_243_0 <= 1'b0;
      shiftRegs_validIn_delay_243_1 <= 1'b0;
      shiftRegs_validIn_delay_244_0 <= 1'b0;
      shiftRegs_validIn_delay_244_1 <= 1'b0;
      shiftRegs_validIn_delay_245_0 <= 1'b0;
      shiftRegs_validIn_delay_245_1 <= 1'b0;
      shiftRegs_validIn_delay_246_0 <= 1'b0;
      shiftRegs_validIn_delay_246_1 <= 1'b0;
      shiftRegs_validIn_delay_247_0 <= 1'b0;
      shiftRegs_validIn_delay_247_1 <= 1'b0;
      shiftRegs_validIn_delay_248_0 <= 1'b0;
      shiftRegs_validIn_delay_248_1 <= 1'b0;
      shiftRegs_validIn_delay_249_0 <= 1'b0;
      shiftRegs_validIn_delay_249_1 <= 1'b0;
      shiftRegs_validIn_delay_250_0 <= 1'b0;
      shiftRegs_validIn_delay_250_1 <= 1'b0;
      shiftRegs_validIn_delay_251_0 <= 1'b0;
      shiftRegs_validIn_delay_251_1 <= 1'b0;
      shiftRegs_validIn_delay_252_0 <= 1'b0;
      shiftRegs_validIn_delay_252_1 <= 1'b0;
      shiftRegs_validIn_delay_253_0 <= 1'b0;
      shiftRegs_validIn_delay_253_1 <= 1'b0;
      shiftRegs_validIn_delay_254_0 <= 1'b0;
      shiftRegs_validIn_delay_254_1 <= 1'b0;
      shiftRegs_validOut_0 <= 1'b0;
      shiftRegs_validOut_1 <= 1'b0;
      shiftRegs_validOut_delay_1_0 <= 1'b0;
      shiftRegs_validOut_delay_1_1 <= 1'b0;
      shiftRegs_validOut_delay_2_0 <= 1'b0;
      shiftRegs_validOut_delay_2_1 <= 1'b0;
      shiftRegs_validOut_delay_3_0 <= 1'b0;
      shiftRegs_validOut_delay_3_1 <= 1'b0;
      shiftRegs_validOut_delay_4_0 <= 1'b0;
      shiftRegs_validOut_delay_4_1 <= 1'b0;
      shiftRegs_validOutFull_0 <= 1'b0;
      shiftRegs_validOutFull_1 <= 1'b0;
      outputValid <= 1'b0;
      flushing_flushCnt_value <= 16'h0;
      flushing_flushCnt_willOverflowIfInc <= 1'b0;
      stage1_NCnt_value <= 32'h0;
      stage1_NCnt_willOverflowIfInc <= 1'b0;
      stage1_GCnt_value <= 4'b0000;
      stage1_GCnt_willOverflowIfInc <= 1'b0;
      stage1_waitReg <= 1'b0;
      stage1_emptyCnt_value <= 9'h0;
      stage1_emptyCnt_willOverflowIfInc <= 1'b0;
      stage1_needAdd1_0 <= 1'b0;
      _zz_stage1_inputValid_0 <= 1'b0;
      _zz_stage1_inputValid_0_1 <= 1'b0;
      _zz_stage1_inputValid_0_2 <= 1'b0;
      _zz_stage1_inputValid_0_3 <= 1'b0;
      _zz_stage1_inputValid_0_4 <= 1'b0;
      stage1_inputValid_0 <= 1'b0;
      _zz_stage1_inputValid_1 <= 1'b0;
      _zz_stage1_inputValid_1_1 <= 1'b0;
      _zz_stage1_inputValid_1_2 <= 1'b0;
      _zz_stage1_inputValid_1_3 <= 1'b0;
      _zz_stage1_inputValid_1_4 <= 1'b0;
      stage1_inputValid_1 <= 1'b0;
      stage2_wCnt_value <= 12'hfff;
      stage2_wCnt_willUnderflowIfDec <= 1'b0;
      stage2_GCnt_value <= 4'b0000;
      stage2_GCnt_willOverflowIfInc <= 1'b0;
      stage2_calCnt_value <= 2'b10;
      stage2_calCnt_willUnderflowIfDec <= 1'b0;
      stage2_waitReg <= 1'b0;
      stage2_waitCnt_value <= 9'h0;
      stage2_waitCnt_willOverflowIfInc <= 1'b0;
      stage3_GCnt_value <= 4'b1001;
      stage3_GCnt_willUnderflowIfDec <= 1'b0;
      stage3_doubleCnt_value <= 5'h0;
      stage3_doubleCnt_willOverflowIfInc <= 1'b0;
      stage3_doubleWaitCnt_value <= 9'h0;
      stage3_doubleWaitCnt_willOverflowIfInc <= 1'b0;
      stage3_addReg <= 1'b0;
      stage3_addWaitCnt_value <= 9'h0;
      stage3_addWaitCnt_willOverflowIfInc <= 1'b0;
      stage3Final_doubleCnt_value <= 4'b0000;
      stage3Final_doubleCnt_willOverflowIfInc <= 1'b0;
      stage3Final_doubleWaitCnt_value <= 9'h0;
      stage3Final_doubleWaitCnt_willOverflowIfInc <= 1'b0;
      stage3Final_addReg <= 1'b0;
      stage3Final_addWaitCnt_value <= 9'h0;
      stage3Final_addWaitCnt_willOverflowIfInc <= 1'b0;
      stage3Final_pAddShr <= 1'b1;
      fsm_stateReg <= fsm_enumDef_flushing;
    end else begin
      if(io_dataIn_valid) begin
        dataInBuffer_validReg <= 1'b1;
      end else begin
        if(dataInBuffer_bufferOut_ready) begin
          dataInBuffer_validReg <= 1'b0;
        end
      end
      shiftRegs_validIn_delay_1_0 <= shiftRegs_validIn_0;
      shiftRegs_validIn_delay_1_1 <= shiftRegs_validIn_1;
      shiftRegs_validIn_delay_2_0 <= shiftRegs_validIn_delay_1_0;
      shiftRegs_validIn_delay_2_1 <= shiftRegs_validIn_delay_1_1;
      shiftRegs_validIn_delay_3_0 <= shiftRegs_validIn_delay_2_0;
      shiftRegs_validIn_delay_3_1 <= shiftRegs_validIn_delay_2_1;
      shiftRegs_validIn_delay_4_0 <= shiftRegs_validIn_delay_3_0;
      shiftRegs_validIn_delay_4_1 <= shiftRegs_validIn_delay_3_1;
      shiftRegs_validIn_delay_5_0 <= shiftRegs_validIn_delay_4_0;
      shiftRegs_validIn_delay_5_1 <= shiftRegs_validIn_delay_4_1;
      shiftRegs_validIn_delay_6_0 <= shiftRegs_validIn_delay_5_0;
      shiftRegs_validIn_delay_6_1 <= shiftRegs_validIn_delay_5_1;
      shiftRegs_validIn_delay_7_0 <= shiftRegs_validIn_delay_6_0;
      shiftRegs_validIn_delay_7_1 <= shiftRegs_validIn_delay_6_1;
      shiftRegs_validIn_delay_8_0 <= shiftRegs_validIn_delay_7_0;
      shiftRegs_validIn_delay_8_1 <= shiftRegs_validIn_delay_7_1;
      shiftRegs_validIn_delay_9_0 <= shiftRegs_validIn_delay_8_0;
      shiftRegs_validIn_delay_9_1 <= shiftRegs_validIn_delay_8_1;
      shiftRegs_validIn_delay_10_0 <= shiftRegs_validIn_delay_9_0;
      shiftRegs_validIn_delay_10_1 <= shiftRegs_validIn_delay_9_1;
      shiftRegs_validIn_delay_11_0 <= shiftRegs_validIn_delay_10_0;
      shiftRegs_validIn_delay_11_1 <= shiftRegs_validIn_delay_10_1;
      shiftRegs_validIn_delay_12_0 <= shiftRegs_validIn_delay_11_0;
      shiftRegs_validIn_delay_12_1 <= shiftRegs_validIn_delay_11_1;
      shiftRegs_validIn_delay_13_0 <= shiftRegs_validIn_delay_12_0;
      shiftRegs_validIn_delay_13_1 <= shiftRegs_validIn_delay_12_1;
      shiftRegs_validIn_delay_14_0 <= shiftRegs_validIn_delay_13_0;
      shiftRegs_validIn_delay_14_1 <= shiftRegs_validIn_delay_13_1;
      shiftRegs_validIn_delay_15_0 <= shiftRegs_validIn_delay_14_0;
      shiftRegs_validIn_delay_15_1 <= shiftRegs_validIn_delay_14_1;
      shiftRegs_validIn_delay_16_0 <= shiftRegs_validIn_delay_15_0;
      shiftRegs_validIn_delay_16_1 <= shiftRegs_validIn_delay_15_1;
      shiftRegs_validIn_delay_17_0 <= shiftRegs_validIn_delay_16_0;
      shiftRegs_validIn_delay_17_1 <= shiftRegs_validIn_delay_16_1;
      shiftRegs_validIn_delay_18_0 <= shiftRegs_validIn_delay_17_0;
      shiftRegs_validIn_delay_18_1 <= shiftRegs_validIn_delay_17_1;
      shiftRegs_validIn_delay_19_0 <= shiftRegs_validIn_delay_18_0;
      shiftRegs_validIn_delay_19_1 <= shiftRegs_validIn_delay_18_1;
      shiftRegs_validIn_delay_20_0 <= shiftRegs_validIn_delay_19_0;
      shiftRegs_validIn_delay_20_1 <= shiftRegs_validIn_delay_19_1;
      shiftRegs_validIn_delay_21_0 <= shiftRegs_validIn_delay_20_0;
      shiftRegs_validIn_delay_21_1 <= shiftRegs_validIn_delay_20_1;
      shiftRegs_validIn_delay_22_0 <= shiftRegs_validIn_delay_21_0;
      shiftRegs_validIn_delay_22_1 <= shiftRegs_validIn_delay_21_1;
      shiftRegs_validIn_delay_23_0 <= shiftRegs_validIn_delay_22_0;
      shiftRegs_validIn_delay_23_1 <= shiftRegs_validIn_delay_22_1;
      shiftRegs_validIn_delay_24_0 <= shiftRegs_validIn_delay_23_0;
      shiftRegs_validIn_delay_24_1 <= shiftRegs_validIn_delay_23_1;
      shiftRegs_validIn_delay_25_0 <= shiftRegs_validIn_delay_24_0;
      shiftRegs_validIn_delay_25_1 <= shiftRegs_validIn_delay_24_1;
      shiftRegs_validIn_delay_26_0 <= shiftRegs_validIn_delay_25_0;
      shiftRegs_validIn_delay_26_1 <= shiftRegs_validIn_delay_25_1;
      shiftRegs_validIn_delay_27_0 <= shiftRegs_validIn_delay_26_0;
      shiftRegs_validIn_delay_27_1 <= shiftRegs_validIn_delay_26_1;
      shiftRegs_validIn_delay_28_0 <= shiftRegs_validIn_delay_27_0;
      shiftRegs_validIn_delay_28_1 <= shiftRegs_validIn_delay_27_1;
      shiftRegs_validIn_delay_29_0 <= shiftRegs_validIn_delay_28_0;
      shiftRegs_validIn_delay_29_1 <= shiftRegs_validIn_delay_28_1;
      shiftRegs_validIn_delay_30_0 <= shiftRegs_validIn_delay_29_0;
      shiftRegs_validIn_delay_30_1 <= shiftRegs_validIn_delay_29_1;
      shiftRegs_validIn_delay_31_0 <= shiftRegs_validIn_delay_30_0;
      shiftRegs_validIn_delay_31_1 <= shiftRegs_validIn_delay_30_1;
      shiftRegs_validIn_delay_32_0 <= shiftRegs_validIn_delay_31_0;
      shiftRegs_validIn_delay_32_1 <= shiftRegs_validIn_delay_31_1;
      shiftRegs_validIn_delay_33_0 <= shiftRegs_validIn_delay_32_0;
      shiftRegs_validIn_delay_33_1 <= shiftRegs_validIn_delay_32_1;
      shiftRegs_validIn_delay_34_0 <= shiftRegs_validIn_delay_33_0;
      shiftRegs_validIn_delay_34_1 <= shiftRegs_validIn_delay_33_1;
      shiftRegs_validIn_delay_35_0 <= shiftRegs_validIn_delay_34_0;
      shiftRegs_validIn_delay_35_1 <= shiftRegs_validIn_delay_34_1;
      shiftRegs_validIn_delay_36_0 <= shiftRegs_validIn_delay_35_0;
      shiftRegs_validIn_delay_36_1 <= shiftRegs_validIn_delay_35_1;
      shiftRegs_validIn_delay_37_0 <= shiftRegs_validIn_delay_36_0;
      shiftRegs_validIn_delay_37_1 <= shiftRegs_validIn_delay_36_1;
      shiftRegs_validIn_delay_38_0 <= shiftRegs_validIn_delay_37_0;
      shiftRegs_validIn_delay_38_1 <= shiftRegs_validIn_delay_37_1;
      shiftRegs_validIn_delay_39_0 <= shiftRegs_validIn_delay_38_0;
      shiftRegs_validIn_delay_39_1 <= shiftRegs_validIn_delay_38_1;
      shiftRegs_validIn_delay_40_0 <= shiftRegs_validIn_delay_39_0;
      shiftRegs_validIn_delay_40_1 <= shiftRegs_validIn_delay_39_1;
      shiftRegs_validIn_delay_41_0 <= shiftRegs_validIn_delay_40_0;
      shiftRegs_validIn_delay_41_1 <= shiftRegs_validIn_delay_40_1;
      shiftRegs_validIn_delay_42_0 <= shiftRegs_validIn_delay_41_0;
      shiftRegs_validIn_delay_42_1 <= shiftRegs_validIn_delay_41_1;
      shiftRegs_validIn_delay_43_0 <= shiftRegs_validIn_delay_42_0;
      shiftRegs_validIn_delay_43_1 <= shiftRegs_validIn_delay_42_1;
      shiftRegs_validIn_delay_44_0 <= shiftRegs_validIn_delay_43_0;
      shiftRegs_validIn_delay_44_1 <= shiftRegs_validIn_delay_43_1;
      shiftRegs_validIn_delay_45_0 <= shiftRegs_validIn_delay_44_0;
      shiftRegs_validIn_delay_45_1 <= shiftRegs_validIn_delay_44_1;
      shiftRegs_validIn_delay_46_0 <= shiftRegs_validIn_delay_45_0;
      shiftRegs_validIn_delay_46_1 <= shiftRegs_validIn_delay_45_1;
      shiftRegs_validIn_delay_47_0 <= shiftRegs_validIn_delay_46_0;
      shiftRegs_validIn_delay_47_1 <= shiftRegs_validIn_delay_46_1;
      shiftRegs_validIn_delay_48_0 <= shiftRegs_validIn_delay_47_0;
      shiftRegs_validIn_delay_48_1 <= shiftRegs_validIn_delay_47_1;
      shiftRegs_validIn_delay_49_0 <= shiftRegs_validIn_delay_48_0;
      shiftRegs_validIn_delay_49_1 <= shiftRegs_validIn_delay_48_1;
      shiftRegs_validIn_delay_50_0 <= shiftRegs_validIn_delay_49_0;
      shiftRegs_validIn_delay_50_1 <= shiftRegs_validIn_delay_49_1;
      shiftRegs_validIn_delay_51_0 <= shiftRegs_validIn_delay_50_0;
      shiftRegs_validIn_delay_51_1 <= shiftRegs_validIn_delay_50_1;
      shiftRegs_validIn_delay_52_0 <= shiftRegs_validIn_delay_51_0;
      shiftRegs_validIn_delay_52_1 <= shiftRegs_validIn_delay_51_1;
      shiftRegs_validIn_delay_53_0 <= shiftRegs_validIn_delay_52_0;
      shiftRegs_validIn_delay_53_1 <= shiftRegs_validIn_delay_52_1;
      shiftRegs_validIn_delay_54_0 <= shiftRegs_validIn_delay_53_0;
      shiftRegs_validIn_delay_54_1 <= shiftRegs_validIn_delay_53_1;
      shiftRegs_validIn_delay_55_0 <= shiftRegs_validIn_delay_54_0;
      shiftRegs_validIn_delay_55_1 <= shiftRegs_validIn_delay_54_1;
      shiftRegs_validIn_delay_56_0 <= shiftRegs_validIn_delay_55_0;
      shiftRegs_validIn_delay_56_1 <= shiftRegs_validIn_delay_55_1;
      shiftRegs_validIn_delay_57_0 <= shiftRegs_validIn_delay_56_0;
      shiftRegs_validIn_delay_57_1 <= shiftRegs_validIn_delay_56_1;
      shiftRegs_validIn_delay_58_0 <= shiftRegs_validIn_delay_57_0;
      shiftRegs_validIn_delay_58_1 <= shiftRegs_validIn_delay_57_1;
      shiftRegs_validIn_delay_59_0 <= shiftRegs_validIn_delay_58_0;
      shiftRegs_validIn_delay_59_1 <= shiftRegs_validIn_delay_58_1;
      shiftRegs_validIn_delay_60_0 <= shiftRegs_validIn_delay_59_0;
      shiftRegs_validIn_delay_60_1 <= shiftRegs_validIn_delay_59_1;
      shiftRegs_validIn_delay_61_0 <= shiftRegs_validIn_delay_60_0;
      shiftRegs_validIn_delay_61_1 <= shiftRegs_validIn_delay_60_1;
      shiftRegs_validIn_delay_62_0 <= shiftRegs_validIn_delay_61_0;
      shiftRegs_validIn_delay_62_1 <= shiftRegs_validIn_delay_61_1;
      shiftRegs_validIn_delay_63_0 <= shiftRegs_validIn_delay_62_0;
      shiftRegs_validIn_delay_63_1 <= shiftRegs_validIn_delay_62_1;
      shiftRegs_validIn_delay_64_0 <= shiftRegs_validIn_delay_63_0;
      shiftRegs_validIn_delay_64_1 <= shiftRegs_validIn_delay_63_1;
      shiftRegs_validIn_delay_65_0 <= shiftRegs_validIn_delay_64_0;
      shiftRegs_validIn_delay_65_1 <= shiftRegs_validIn_delay_64_1;
      shiftRegs_validIn_delay_66_0 <= shiftRegs_validIn_delay_65_0;
      shiftRegs_validIn_delay_66_1 <= shiftRegs_validIn_delay_65_1;
      shiftRegs_validIn_delay_67_0 <= shiftRegs_validIn_delay_66_0;
      shiftRegs_validIn_delay_67_1 <= shiftRegs_validIn_delay_66_1;
      shiftRegs_validIn_delay_68_0 <= shiftRegs_validIn_delay_67_0;
      shiftRegs_validIn_delay_68_1 <= shiftRegs_validIn_delay_67_1;
      shiftRegs_validIn_delay_69_0 <= shiftRegs_validIn_delay_68_0;
      shiftRegs_validIn_delay_69_1 <= shiftRegs_validIn_delay_68_1;
      shiftRegs_validIn_delay_70_0 <= shiftRegs_validIn_delay_69_0;
      shiftRegs_validIn_delay_70_1 <= shiftRegs_validIn_delay_69_1;
      shiftRegs_validIn_delay_71_0 <= shiftRegs_validIn_delay_70_0;
      shiftRegs_validIn_delay_71_1 <= shiftRegs_validIn_delay_70_1;
      shiftRegs_validIn_delay_72_0 <= shiftRegs_validIn_delay_71_0;
      shiftRegs_validIn_delay_72_1 <= shiftRegs_validIn_delay_71_1;
      shiftRegs_validIn_delay_73_0 <= shiftRegs_validIn_delay_72_0;
      shiftRegs_validIn_delay_73_1 <= shiftRegs_validIn_delay_72_1;
      shiftRegs_validIn_delay_74_0 <= shiftRegs_validIn_delay_73_0;
      shiftRegs_validIn_delay_74_1 <= shiftRegs_validIn_delay_73_1;
      shiftRegs_validIn_delay_75_0 <= shiftRegs_validIn_delay_74_0;
      shiftRegs_validIn_delay_75_1 <= shiftRegs_validIn_delay_74_1;
      shiftRegs_validIn_delay_76_0 <= shiftRegs_validIn_delay_75_0;
      shiftRegs_validIn_delay_76_1 <= shiftRegs_validIn_delay_75_1;
      shiftRegs_validIn_delay_77_0 <= shiftRegs_validIn_delay_76_0;
      shiftRegs_validIn_delay_77_1 <= shiftRegs_validIn_delay_76_1;
      shiftRegs_validIn_delay_78_0 <= shiftRegs_validIn_delay_77_0;
      shiftRegs_validIn_delay_78_1 <= shiftRegs_validIn_delay_77_1;
      shiftRegs_validIn_delay_79_0 <= shiftRegs_validIn_delay_78_0;
      shiftRegs_validIn_delay_79_1 <= shiftRegs_validIn_delay_78_1;
      shiftRegs_validIn_delay_80_0 <= shiftRegs_validIn_delay_79_0;
      shiftRegs_validIn_delay_80_1 <= shiftRegs_validIn_delay_79_1;
      shiftRegs_validIn_delay_81_0 <= shiftRegs_validIn_delay_80_0;
      shiftRegs_validIn_delay_81_1 <= shiftRegs_validIn_delay_80_1;
      shiftRegs_validIn_delay_82_0 <= shiftRegs_validIn_delay_81_0;
      shiftRegs_validIn_delay_82_1 <= shiftRegs_validIn_delay_81_1;
      shiftRegs_validIn_delay_83_0 <= shiftRegs_validIn_delay_82_0;
      shiftRegs_validIn_delay_83_1 <= shiftRegs_validIn_delay_82_1;
      shiftRegs_validIn_delay_84_0 <= shiftRegs_validIn_delay_83_0;
      shiftRegs_validIn_delay_84_1 <= shiftRegs_validIn_delay_83_1;
      shiftRegs_validIn_delay_85_0 <= shiftRegs_validIn_delay_84_0;
      shiftRegs_validIn_delay_85_1 <= shiftRegs_validIn_delay_84_1;
      shiftRegs_validIn_delay_86_0 <= shiftRegs_validIn_delay_85_0;
      shiftRegs_validIn_delay_86_1 <= shiftRegs_validIn_delay_85_1;
      shiftRegs_validIn_delay_87_0 <= shiftRegs_validIn_delay_86_0;
      shiftRegs_validIn_delay_87_1 <= shiftRegs_validIn_delay_86_1;
      shiftRegs_validIn_delay_88_0 <= shiftRegs_validIn_delay_87_0;
      shiftRegs_validIn_delay_88_1 <= shiftRegs_validIn_delay_87_1;
      shiftRegs_validIn_delay_89_0 <= shiftRegs_validIn_delay_88_0;
      shiftRegs_validIn_delay_89_1 <= shiftRegs_validIn_delay_88_1;
      shiftRegs_validIn_delay_90_0 <= shiftRegs_validIn_delay_89_0;
      shiftRegs_validIn_delay_90_1 <= shiftRegs_validIn_delay_89_1;
      shiftRegs_validIn_delay_91_0 <= shiftRegs_validIn_delay_90_0;
      shiftRegs_validIn_delay_91_1 <= shiftRegs_validIn_delay_90_1;
      shiftRegs_validIn_delay_92_0 <= shiftRegs_validIn_delay_91_0;
      shiftRegs_validIn_delay_92_1 <= shiftRegs_validIn_delay_91_1;
      shiftRegs_validIn_delay_93_0 <= shiftRegs_validIn_delay_92_0;
      shiftRegs_validIn_delay_93_1 <= shiftRegs_validIn_delay_92_1;
      shiftRegs_validIn_delay_94_0 <= shiftRegs_validIn_delay_93_0;
      shiftRegs_validIn_delay_94_1 <= shiftRegs_validIn_delay_93_1;
      shiftRegs_validIn_delay_95_0 <= shiftRegs_validIn_delay_94_0;
      shiftRegs_validIn_delay_95_1 <= shiftRegs_validIn_delay_94_1;
      shiftRegs_validIn_delay_96_0 <= shiftRegs_validIn_delay_95_0;
      shiftRegs_validIn_delay_96_1 <= shiftRegs_validIn_delay_95_1;
      shiftRegs_validIn_delay_97_0 <= shiftRegs_validIn_delay_96_0;
      shiftRegs_validIn_delay_97_1 <= shiftRegs_validIn_delay_96_1;
      shiftRegs_validIn_delay_98_0 <= shiftRegs_validIn_delay_97_0;
      shiftRegs_validIn_delay_98_1 <= shiftRegs_validIn_delay_97_1;
      shiftRegs_validIn_delay_99_0 <= shiftRegs_validIn_delay_98_0;
      shiftRegs_validIn_delay_99_1 <= shiftRegs_validIn_delay_98_1;
      shiftRegs_validIn_delay_100_0 <= shiftRegs_validIn_delay_99_0;
      shiftRegs_validIn_delay_100_1 <= shiftRegs_validIn_delay_99_1;
      shiftRegs_validIn_delay_101_0 <= shiftRegs_validIn_delay_100_0;
      shiftRegs_validIn_delay_101_1 <= shiftRegs_validIn_delay_100_1;
      shiftRegs_validIn_delay_102_0 <= shiftRegs_validIn_delay_101_0;
      shiftRegs_validIn_delay_102_1 <= shiftRegs_validIn_delay_101_1;
      shiftRegs_validIn_delay_103_0 <= shiftRegs_validIn_delay_102_0;
      shiftRegs_validIn_delay_103_1 <= shiftRegs_validIn_delay_102_1;
      shiftRegs_validIn_delay_104_0 <= shiftRegs_validIn_delay_103_0;
      shiftRegs_validIn_delay_104_1 <= shiftRegs_validIn_delay_103_1;
      shiftRegs_validIn_delay_105_0 <= shiftRegs_validIn_delay_104_0;
      shiftRegs_validIn_delay_105_1 <= shiftRegs_validIn_delay_104_1;
      shiftRegs_validIn_delay_106_0 <= shiftRegs_validIn_delay_105_0;
      shiftRegs_validIn_delay_106_1 <= shiftRegs_validIn_delay_105_1;
      shiftRegs_validIn_delay_107_0 <= shiftRegs_validIn_delay_106_0;
      shiftRegs_validIn_delay_107_1 <= shiftRegs_validIn_delay_106_1;
      shiftRegs_validIn_delay_108_0 <= shiftRegs_validIn_delay_107_0;
      shiftRegs_validIn_delay_108_1 <= shiftRegs_validIn_delay_107_1;
      shiftRegs_validIn_delay_109_0 <= shiftRegs_validIn_delay_108_0;
      shiftRegs_validIn_delay_109_1 <= shiftRegs_validIn_delay_108_1;
      shiftRegs_validIn_delay_110_0 <= shiftRegs_validIn_delay_109_0;
      shiftRegs_validIn_delay_110_1 <= shiftRegs_validIn_delay_109_1;
      shiftRegs_validIn_delay_111_0 <= shiftRegs_validIn_delay_110_0;
      shiftRegs_validIn_delay_111_1 <= shiftRegs_validIn_delay_110_1;
      shiftRegs_validIn_delay_112_0 <= shiftRegs_validIn_delay_111_0;
      shiftRegs_validIn_delay_112_1 <= shiftRegs_validIn_delay_111_1;
      shiftRegs_validIn_delay_113_0 <= shiftRegs_validIn_delay_112_0;
      shiftRegs_validIn_delay_113_1 <= shiftRegs_validIn_delay_112_1;
      shiftRegs_validIn_delay_114_0 <= shiftRegs_validIn_delay_113_0;
      shiftRegs_validIn_delay_114_1 <= shiftRegs_validIn_delay_113_1;
      shiftRegs_validIn_delay_115_0 <= shiftRegs_validIn_delay_114_0;
      shiftRegs_validIn_delay_115_1 <= shiftRegs_validIn_delay_114_1;
      shiftRegs_validIn_delay_116_0 <= shiftRegs_validIn_delay_115_0;
      shiftRegs_validIn_delay_116_1 <= shiftRegs_validIn_delay_115_1;
      shiftRegs_validIn_delay_117_0 <= shiftRegs_validIn_delay_116_0;
      shiftRegs_validIn_delay_117_1 <= shiftRegs_validIn_delay_116_1;
      shiftRegs_validIn_delay_118_0 <= shiftRegs_validIn_delay_117_0;
      shiftRegs_validIn_delay_118_1 <= shiftRegs_validIn_delay_117_1;
      shiftRegs_validIn_delay_119_0 <= shiftRegs_validIn_delay_118_0;
      shiftRegs_validIn_delay_119_1 <= shiftRegs_validIn_delay_118_1;
      shiftRegs_validIn_delay_120_0 <= shiftRegs_validIn_delay_119_0;
      shiftRegs_validIn_delay_120_1 <= shiftRegs_validIn_delay_119_1;
      shiftRegs_validIn_delay_121_0 <= shiftRegs_validIn_delay_120_0;
      shiftRegs_validIn_delay_121_1 <= shiftRegs_validIn_delay_120_1;
      shiftRegs_validIn_delay_122_0 <= shiftRegs_validIn_delay_121_0;
      shiftRegs_validIn_delay_122_1 <= shiftRegs_validIn_delay_121_1;
      shiftRegs_validIn_delay_123_0 <= shiftRegs_validIn_delay_122_0;
      shiftRegs_validIn_delay_123_1 <= shiftRegs_validIn_delay_122_1;
      shiftRegs_validIn_delay_124_0 <= shiftRegs_validIn_delay_123_0;
      shiftRegs_validIn_delay_124_1 <= shiftRegs_validIn_delay_123_1;
      shiftRegs_validIn_delay_125_0 <= shiftRegs_validIn_delay_124_0;
      shiftRegs_validIn_delay_125_1 <= shiftRegs_validIn_delay_124_1;
      shiftRegs_validIn_delay_126_0 <= shiftRegs_validIn_delay_125_0;
      shiftRegs_validIn_delay_126_1 <= shiftRegs_validIn_delay_125_1;
      shiftRegs_validIn_delay_127_0 <= shiftRegs_validIn_delay_126_0;
      shiftRegs_validIn_delay_127_1 <= shiftRegs_validIn_delay_126_1;
      shiftRegs_validIn_delay_128_0 <= shiftRegs_validIn_delay_127_0;
      shiftRegs_validIn_delay_128_1 <= shiftRegs_validIn_delay_127_1;
      shiftRegs_validIn_delay_129_0 <= shiftRegs_validIn_delay_128_0;
      shiftRegs_validIn_delay_129_1 <= shiftRegs_validIn_delay_128_1;
      shiftRegs_validIn_delay_130_0 <= shiftRegs_validIn_delay_129_0;
      shiftRegs_validIn_delay_130_1 <= shiftRegs_validIn_delay_129_1;
      shiftRegs_validIn_delay_131_0 <= shiftRegs_validIn_delay_130_0;
      shiftRegs_validIn_delay_131_1 <= shiftRegs_validIn_delay_130_1;
      shiftRegs_validIn_delay_132_0 <= shiftRegs_validIn_delay_131_0;
      shiftRegs_validIn_delay_132_1 <= shiftRegs_validIn_delay_131_1;
      shiftRegs_validIn_delay_133_0 <= shiftRegs_validIn_delay_132_0;
      shiftRegs_validIn_delay_133_1 <= shiftRegs_validIn_delay_132_1;
      shiftRegs_validIn_delay_134_0 <= shiftRegs_validIn_delay_133_0;
      shiftRegs_validIn_delay_134_1 <= shiftRegs_validIn_delay_133_1;
      shiftRegs_validIn_delay_135_0 <= shiftRegs_validIn_delay_134_0;
      shiftRegs_validIn_delay_135_1 <= shiftRegs_validIn_delay_134_1;
      shiftRegs_validIn_delay_136_0 <= shiftRegs_validIn_delay_135_0;
      shiftRegs_validIn_delay_136_1 <= shiftRegs_validIn_delay_135_1;
      shiftRegs_validIn_delay_137_0 <= shiftRegs_validIn_delay_136_0;
      shiftRegs_validIn_delay_137_1 <= shiftRegs_validIn_delay_136_1;
      shiftRegs_validIn_delay_138_0 <= shiftRegs_validIn_delay_137_0;
      shiftRegs_validIn_delay_138_1 <= shiftRegs_validIn_delay_137_1;
      shiftRegs_validIn_delay_139_0 <= shiftRegs_validIn_delay_138_0;
      shiftRegs_validIn_delay_139_1 <= shiftRegs_validIn_delay_138_1;
      shiftRegs_validIn_delay_140_0 <= shiftRegs_validIn_delay_139_0;
      shiftRegs_validIn_delay_140_1 <= shiftRegs_validIn_delay_139_1;
      shiftRegs_validIn_delay_141_0 <= shiftRegs_validIn_delay_140_0;
      shiftRegs_validIn_delay_141_1 <= shiftRegs_validIn_delay_140_1;
      shiftRegs_validIn_delay_142_0 <= shiftRegs_validIn_delay_141_0;
      shiftRegs_validIn_delay_142_1 <= shiftRegs_validIn_delay_141_1;
      shiftRegs_validIn_delay_143_0 <= shiftRegs_validIn_delay_142_0;
      shiftRegs_validIn_delay_143_1 <= shiftRegs_validIn_delay_142_1;
      shiftRegs_validIn_delay_144_0 <= shiftRegs_validIn_delay_143_0;
      shiftRegs_validIn_delay_144_1 <= shiftRegs_validIn_delay_143_1;
      shiftRegs_validIn_delay_145_0 <= shiftRegs_validIn_delay_144_0;
      shiftRegs_validIn_delay_145_1 <= shiftRegs_validIn_delay_144_1;
      shiftRegs_validIn_delay_146_0 <= shiftRegs_validIn_delay_145_0;
      shiftRegs_validIn_delay_146_1 <= shiftRegs_validIn_delay_145_1;
      shiftRegs_validIn_delay_147_0 <= shiftRegs_validIn_delay_146_0;
      shiftRegs_validIn_delay_147_1 <= shiftRegs_validIn_delay_146_1;
      shiftRegs_validIn_delay_148_0 <= shiftRegs_validIn_delay_147_0;
      shiftRegs_validIn_delay_148_1 <= shiftRegs_validIn_delay_147_1;
      shiftRegs_validIn_delay_149_0 <= shiftRegs_validIn_delay_148_0;
      shiftRegs_validIn_delay_149_1 <= shiftRegs_validIn_delay_148_1;
      shiftRegs_validIn_delay_150_0 <= shiftRegs_validIn_delay_149_0;
      shiftRegs_validIn_delay_150_1 <= shiftRegs_validIn_delay_149_1;
      shiftRegs_validIn_delay_151_0 <= shiftRegs_validIn_delay_150_0;
      shiftRegs_validIn_delay_151_1 <= shiftRegs_validIn_delay_150_1;
      shiftRegs_validIn_delay_152_0 <= shiftRegs_validIn_delay_151_0;
      shiftRegs_validIn_delay_152_1 <= shiftRegs_validIn_delay_151_1;
      shiftRegs_validIn_delay_153_0 <= shiftRegs_validIn_delay_152_0;
      shiftRegs_validIn_delay_153_1 <= shiftRegs_validIn_delay_152_1;
      shiftRegs_validIn_delay_154_0 <= shiftRegs_validIn_delay_153_0;
      shiftRegs_validIn_delay_154_1 <= shiftRegs_validIn_delay_153_1;
      shiftRegs_validIn_delay_155_0 <= shiftRegs_validIn_delay_154_0;
      shiftRegs_validIn_delay_155_1 <= shiftRegs_validIn_delay_154_1;
      shiftRegs_validIn_delay_156_0 <= shiftRegs_validIn_delay_155_0;
      shiftRegs_validIn_delay_156_1 <= shiftRegs_validIn_delay_155_1;
      shiftRegs_validIn_delay_157_0 <= shiftRegs_validIn_delay_156_0;
      shiftRegs_validIn_delay_157_1 <= shiftRegs_validIn_delay_156_1;
      shiftRegs_validIn_delay_158_0 <= shiftRegs_validIn_delay_157_0;
      shiftRegs_validIn_delay_158_1 <= shiftRegs_validIn_delay_157_1;
      shiftRegs_validIn_delay_159_0 <= shiftRegs_validIn_delay_158_0;
      shiftRegs_validIn_delay_159_1 <= shiftRegs_validIn_delay_158_1;
      shiftRegs_validIn_delay_160_0 <= shiftRegs_validIn_delay_159_0;
      shiftRegs_validIn_delay_160_1 <= shiftRegs_validIn_delay_159_1;
      shiftRegs_validIn_delay_161_0 <= shiftRegs_validIn_delay_160_0;
      shiftRegs_validIn_delay_161_1 <= shiftRegs_validIn_delay_160_1;
      shiftRegs_validIn_delay_162_0 <= shiftRegs_validIn_delay_161_0;
      shiftRegs_validIn_delay_162_1 <= shiftRegs_validIn_delay_161_1;
      shiftRegs_validIn_delay_163_0 <= shiftRegs_validIn_delay_162_0;
      shiftRegs_validIn_delay_163_1 <= shiftRegs_validIn_delay_162_1;
      shiftRegs_validIn_delay_164_0 <= shiftRegs_validIn_delay_163_0;
      shiftRegs_validIn_delay_164_1 <= shiftRegs_validIn_delay_163_1;
      shiftRegs_validIn_delay_165_0 <= shiftRegs_validIn_delay_164_0;
      shiftRegs_validIn_delay_165_1 <= shiftRegs_validIn_delay_164_1;
      shiftRegs_validIn_delay_166_0 <= shiftRegs_validIn_delay_165_0;
      shiftRegs_validIn_delay_166_1 <= shiftRegs_validIn_delay_165_1;
      shiftRegs_validIn_delay_167_0 <= shiftRegs_validIn_delay_166_0;
      shiftRegs_validIn_delay_167_1 <= shiftRegs_validIn_delay_166_1;
      shiftRegs_validIn_delay_168_0 <= shiftRegs_validIn_delay_167_0;
      shiftRegs_validIn_delay_168_1 <= shiftRegs_validIn_delay_167_1;
      shiftRegs_validIn_delay_169_0 <= shiftRegs_validIn_delay_168_0;
      shiftRegs_validIn_delay_169_1 <= shiftRegs_validIn_delay_168_1;
      shiftRegs_validIn_delay_170_0 <= shiftRegs_validIn_delay_169_0;
      shiftRegs_validIn_delay_170_1 <= shiftRegs_validIn_delay_169_1;
      shiftRegs_validIn_delay_171_0 <= shiftRegs_validIn_delay_170_0;
      shiftRegs_validIn_delay_171_1 <= shiftRegs_validIn_delay_170_1;
      shiftRegs_validIn_delay_172_0 <= shiftRegs_validIn_delay_171_0;
      shiftRegs_validIn_delay_172_1 <= shiftRegs_validIn_delay_171_1;
      shiftRegs_validIn_delay_173_0 <= shiftRegs_validIn_delay_172_0;
      shiftRegs_validIn_delay_173_1 <= shiftRegs_validIn_delay_172_1;
      shiftRegs_validIn_delay_174_0 <= shiftRegs_validIn_delay_173_0;
      shiftRegs_validIn_delay_174_1 <= shiftRegs_validIn_delay_173_1;
      shiftRegs_validIn_delay_175_0 <= shiftRegs_validIn_delay_174_0;
      shiftRegs_validIn_delay_175_1 <= shiftRegs_validIn_delay_174_1;
      shiftRegs_validIn_delay_176_0 <= shiftRegs_validIn_delay_175_0;
      shiftRegs_validIn_delay_176_1 <= shiftRegs_validIn_delay_175_1;
      shiftRegs_validIn_delay_177_0 <= shiftRegs_validIn_delay_176_0;
      shiftRegs_validIn_delay_177_1 <= shiftRegs_validIn_delay_176_1;
      shiftRegs_validIn_delay_178_0 <= shiftRegs_validIn_delay_177_0;
      shiftRegs_validIn_delay_178_1 <= shiftRegs_validIn_delay_177_1;
      shiftRegs_validIn_delay_179_0 <= shiftRegs_validIn_delay_178_0;
      shiftRegs_validIn_delay_179_1 <= shiftRegs_validIn_delay_178_1;
      shiftRegs_validIn_delay_180_0 <= shiftRegs_validIn_delay_179_0;
      shiftRegs_validIn_delay_180_1 <= shiftRegs_validIn_delay_179_1;
      shiftRegs_validIn_delay_181_0 <= shiftRegs_validIn_delay_180_0;
      shiftRegs_validIn_delay_181_1 <= shiftRegs_validIn_delay_180_1;
      shiftRegs_validIn_delay_182_0 <= shiftRegs_validIn_delay_181_0;
      shiftRegs_validIn_delay_182_1 <= shiftRegs_validIn_delay_181_1;
      shiftRegs_validIn_delay_183_0 <= shiftRegs_validIn_delay_182_0;
      shiftRegs_validIn_delay_183_1 <= shiftRegs_validIn_delay_182_1;
      shiftRegs_validIn_delay_184_0 <= shiftRegs_validIn_delay_183_0;
      shiftRegs_validIn_delay_184_1 <= shiftRegs_validIn_delay_183_1;
      shiftRegs_validIn_delay_185_0 <= shiftRegs_validIn_delay_184_0;
      shiftRegs_validIn_delay_185_1 <= shiftRegs_validIn_delay_184_1;
      shiftRegs_validIn_delay_186_0 <= shiftRegs_validIn_delay_185_0;
      shiftRegs_validIn_delay_186_1 <= shiftRegs_validIn_delay_185_1;
      shiftRegs_validIn_delay_187_0 <= shiftRegs_validIn_delay_186_0;
      shiftRegs_validIn_delay_187_1 <= shiftRegs_validIn_delay_186_1;
      shiftRegs_validIn_delay_188_0 <= shiftRegs_validIn_delay_187_0;
      shiftRegs_validIn_delay_188_1 <= shiftRegs_validIn_delay_187_1;
      shiftRegs_validIn_delay_189_0 <= shiftRegs_validIn_delay_188_0;
      shiftRegs_validIn_delay_189_1 <= shiftRegs_validIn_delay_188_1;
      shiftRegs_validIn_delay_190_0 <= shiftRegs_validIn_delay_189_0;
      shiftRegs_validIn_delay_190_1 <= shiftRegs_validIn_delay_189_1;
      shiftRegs_validIn_delay_191_0 <= shiftRegs_validIn_delay_190_0;
      shiftRegs_validIn_delay_191_1 <= shiftRegs_validIn_delay_190_1;
      shiftRegs_validIn_delay_192_0 <= shiftRegs_validIn_delay_191_0;
      shiftRegs_validIn_delay_192_1 <= shiftRegs_validIn_delay_191_1;
      shiftRegs_validIn_delay_193_0 <= shiftRegs_validIn_delay_192_0;
      shiftRegs_validIn_delay_193_1 <= shiftRegs_validIn_delay_192_1;
      shiftRegs_validIn_delay_194_0 <= shiftRegs_validIn_delay_193_0;
      shiftRegs_validIn_delay_194_1 <= shiftRegs_validIn_delay_193_1;
      shiftRegs_validIn_delay_195_0 <= shiftRegs_validIn_delay_194_0;
      shiftRegs_validIn_delay_195_1 <= shiftRegs_validIn_delay_194_1;
      shiftRegs_validIn_delay_196_0 <= shiftRegs_validIn_delay_195_0;
      shiftRegs_validIn_delay_196_1 <= shiftRegs_validIn_delay_195_1;
      shiftRegs_validIn_delay_197_0 <= shiftRegs_validIn_delay_196_0;
      shiftRegs_validIn_delay_197_1 <= shiftRegs_validIn_delay_196_1;
      shiftRegs_validIn_delay_198_0 <= shiftRegs_validIn_delay_197_0;
      shiftRegs_validIn_delay_198_1 <= shiftRegs_validIn_delay_197_1;
      shiftRegs_validIn_delay_199_0 <= shiftRegs_validIn_delay_198_0;
      shiftRegs_validIn_delay_199_1 <= shiftRegs_validIn_delay_198_1;
      shiftRegs_validIn_delay_200_0 <= shiftRegs_validIn_delay_199_0;
      shiftRegs_validIn_delay_200_1 <= shiftRegs_validIn_delay_199_1;
      shiftRegs_validIn_delay_201_0 <= shiftRegs_validIn_delay_200_0;
      shiftRegs_validIn_delay_201_1 <= shiftRegs_validIn_delay_200_1;
      shiftRegs_validIn_delay_202_0 <= shiftRegs_validIn_delay_201_0;
      shiftRegs_validIn_delay_202_1 <= shiftRegs_validIn_delay_201_1;
      shiftRegs_validIn_delay_203_0 <= shiftRegs_validIn_delay_202_0;
      shiftRegs_validIn_delay_203_1 <= shiftRegs_validIn_delay_202_1;
      shiftRegs_validIn_delay_204_0 <= shiftRegs_validIn_delay_203_0;
      shiftRegs_validIn_delay_204_1 <= shiftRegs_validIn_delay_203_1;
      shiftRegs_validIn_delay_205_0 <= shiftRegs_validIn_delay_204_0;
      shiftRegs_validIn_delay_205_1 <= shiftRegs_validIn_delay_204_1;
      shiftRegs_validIn_delay_206_0 <= shiftRegs_validIn_delay_205_0;
      shiftRegs_validIn_delay_206_1 <= shiftRegs_validIn_delay_205_1;
      shiftRegs_validIn_delay_207_0 <= shiftRegs_validIn_delay_206_0;
      shiftRegs_validIn_delay_207_1 <= shiftRegs_validIn_delay_206_1;
      shiftRegs_validIn_delay_208_0 <= shiftRegs_validIn_delay_207_0;
      shiftRegs_validIn_delay_208_1 <= shiftRegs_validIn_delay_207_1;
      shiftRegs_validIn_delay_209_0 <= shiftRegs_validIn_delay_208_0;
      shiftRegs_validIn_delay_209_1 <= shiftRegs_validIn_delay_208_1;
      shiftRegs_validIn_delay_210_0 <= shiftRegs_validIn_delay_209_0;
      shiftRegs_validIn_delay_210_1 <= shiftRegs_validIn_delay_209_1;
      shiftRegs_validIn_delay_211_0 <= shiftRegs_validIn_delay_210_0;
      shiftRegs_validIn_delay_211_1 <= shiftRegs_validIn_delay_210_1;
      shiftRegs_validIn_delay_212_0 <= shiftRegs_validIn_delay_211_0;
      shiftRegs_validIn_delay_212_1 <= shiftRegs_validIn_delay_211_1;
      shiftRegs_validIn_delay_213_0 <= shiftRegs_validIn_delay_212_0;
      shiftRegs_validIn_delay_213_1 <= shiftRegs_validIn_delay_212_1;
      shiftRegs_validIn_delay_214_0 <= shiftRegs_validIn_delay_213_0;
      shiftRegs_validIn_delay_214_1 <= shiftRegs_validIn_delay_213_1;
      shiftRegs_validIn_delay_215_0 <= shiftRegs_validIn_delay_214_0;
      shiftRegs_validIn_delay_215_1 <= shiftRegs_validIn_delay_214_1;
      shiftRegs_validIn_delay_216_0 <= shiftRegs_validIn_delay_215_0;
      shiftRegs_validIn_delay_216_1 <= shiftRegs_validIn_delay_215_1;
      shiftRegs_validIn_delay_217_0 <= shiftRegs_validIn_delay_216_0;
      shiftRegs_validIn_delay_217_1 <= shiftRegs_validIn_delay_216_1;
      shiftRegs_validIn_delay_218_0 <= shiftRegs_validIn_delay_217_0;
      shiftRegs_validIn_delay_218_1 <= shiftRegs_validIn_delay_217_1;
      shiftRegs_validIn_delay_219_0 <= shiftRegs_validIn_delay_218_0;
      shiftRegs_validIn_delay_219_1 <= shiftRegs_validIn_delay_218_1;
      shiftRegs_validIn_delay_220_0 <= shiftRegs_validIn_delay_219_0;
      shiftRegs_validIn_delay_220_1 <= shiftRegs_validIn_delay_219_1;
      shiftRegs_validIn_delay_221_0 <= shiftRegs_validIn_delay_220_0;
      shiftRegs_validIn_delay_221_1 <= shiftRegs_validIn_delay_220_1;
      shiftRegs_validIn_delay_222_0 <= shiftRegs_validIn_delay_221_0;
      shiftRegs_validIn_delay_222_1 <= shiftRegs_validIn_delay_221_1;
      shiftRegs_validIn_delay_223_0 <= shiftRegs_validIn_delay_222_0;
      shiftRegs_validIn_delay_223_1 <= shiftRegs_validIn_delay_222_1;
      shiftRegs_validIn_delay_224_0 <= shiftRegs_validIn_delay_223_0;
      shiftRegs_validIn_delay_224_1 <= shiftRegs_validIn_delay_223_1;
      shiftRegs_validIn_delay_225_0 <= shiftRegs_validIn_delay_224_0;
      shiftRegs_validIn_delay_225_1 <= shiftRegs_validIn_delay_224_1;
      shiftRegs_validIn_delay_226_0 <= shiftRegs_validIn_delay_225_0;
      shiftRegs_validIn_delay_226_1 <= shiftRegs_validIn_delay_225_1;
      shiftRegs_validIn_delay_227_0 <= shiftRegs_validIn_delay_226_0;
      shiftRegs_validIn_delay_227_1 <= shiftRegs_validIn_delay_226_1;
      shiftRegs_validIn_delay_228_0 <= shiftRegs_validIn_delay_227_0;
      shiftRegs_validIn_delay_228_1 <= shiftRegs_validIn_delay_227_1;
      shiftRegs_validIn_delay_229_0 <= shiftRegs_validIn_delay_228_0;
      shiftRegs_validIn_delay_229_1 <= shiftRegs_validIn_delay_228_1;
      shiftRegs_validIn_delay_230_0 <= shiftRegs_validIn_delay_229_0;
      shiftRegs_validIn_delay_230_1 <= shiftRegs_validIn_delay_229_1;
      shiftRegs_validIn_delay_231_0 <= shiftRegs_validIn_delay_230_0;
      shiftRegs_validIn_delay_231_1 <= shiftRegs_validIn_delay_230_1;
      shiftRegs_validIn_delay_232_0 <= shiftRegs_validIn_delay_231_0;
      shiftRegs_validIn_delay_232_1 <= shiftRegs_validIn_delay_231_1;
      shiftRegs_validIn_delay_233_0 <= shiftRegs_validIn_delay_232_0;
      shiftRegs_validIn_delay_233_1 <= shiftRegs_validIn_delay_232_1;
      shiftRegs_validIn_delay_234_0 <= shiftRegs_validIn_delay_233_0;
      shiftRegs_validIn_delay_234_1 <= shiftRegs_validIn_delay_233_1;
      shiftRegs_validIn_delay_235_0 <= shiftRegs_validIn_delay_234_0;
      shiftRegs_validIn_delay_235_1 <= shiftRegs_validIn_delay_234_1;
      shiftRegs_validIn_delay_236_0 <= shiftRegs_validIn_delay_235_0;
      shiftRegs_validIn_delay_236_1 <= shiftRegs_validIn_delay_235_1;
      shiftRegs_validIn_delay_237_0 <= shiftRegs_validIn_delay_236_0;
      shiftRegs_validIn_delay_237_1 <= shiftRegs_validIn_delay_236_1;
      shiftRegs_validIn_delay_238_0 <= shiftRegs_validIn_delay_237_0;
      shiftRegs_validIn_delay_238_1 <= shiftRegs_validIn_delay_237_1;
      shiftRegs_validIn_delay_239_0 <= shiftRegs_validIn_delay_238_0;
      shiftRegs_validIn_delay_239_1 <= shiftRegs_validIn_delay_238_1;
      shiftRegs_validIn_delay_240_0 <= shiftRegs_validIn_delay_239_0;
      shiftRegs_validIn_delay_240_1 <= shiftRegs_validIn_delay_239_1;
      shiftRegs_validIn_delay_241_0 <= shiftRegs_validIn_delay_240_0;
      shiftRegs_validIn_delay_241_1 <= shiftRegs_validIn_delay_240_1;
      shiftRegs_validIn_delay_242_0 <= shiftRegs_validIn_delay_241_0;
      shiftRegs_validIn_delay_242_1 <= shiftRegs_validIn_delay_241_1;
      shiftRegs_validIn_delay_243_0 <= shiftRegs_validIn_delay_242_0;
      shiftRegs_validIn_delay_243_1 <= shiftRegs_validIn_delay_242_1;
      shiftRegs_validIn_delay_244_0 <= shiftRegs_validIn_delay_243_0;
      shiftRegs_validIn_delay_244_1 <= shiftRegs_validIn_delay_243_1;
      shiftRegs_validIn_delay_245_0 <= shiftRegs_validIn_delay_244_0;
      shiftRegs_validIn_delay_245_1 <= shiftRegs_validIn_delay_244_1;
      shiftRegs_validIn_delay_246_0 <= shiftRegs_validIn_delay_245_0;
      shiftRegs_validIn_delay_246_1 <= shiftRegs_validIn_delay_245_1;
      shiftRegs_validIn_delay_247_0 <= shiftRegs_validIn_delay_246_0;
      shiftRegs_validIn_delay_247_1 <= shiftRegs_validIn_delay_246_1;
      shiftRegs_validIn_delay_248_0 <= shiftRegs_validIn_delay_247_0;
      shiftRegs_validIn_delay_248_1 <= shiftRegs_validIn_delay_247_1;
      shiftRegs_validIn_delay_249_0 <= shiftRegs_validIn_delay_248_0;
      shiftRegs_validIn_delay_249_1 <= shiftRegs_validIn_delay_248_1;
      shiftRegs_validIn_delay_250_0 <= shiftRegs_validIn_delay_249_0;
      shiftRegs_validIn_delay_250_1 <= shiftRegs_validIn_delay_249_1;
      shiftRegs_validIn_delay_251_0 <= shiftRegs_validIn_delay_250_0;
      shiftRegs_validIn_delay_251_1 <= shiftRegs_validIn_delay_250_1;
      shiftRegs_validIn_delay_252_0 <= shiftRegs_validIn_delay_251_0;
      shiftRegs_validIn_delay_252_1 <= shiftRegs_validIn_delay_251_1;
      shiftRegs_validIn_delay_253_0 <= shiftRegs_validIn_delay_252_0;
      shiftRegs_validIn_delay_253_1 <= shiftRegs_validIn_delay_252_1;
      shiftRegs_validIn_delay_254_0 <= shiftRegs_validIn_delay_253_0;
      shiftRegs_validIn_delay_254_1 <= shiftRegs_validIn_delay_253_1;
      shiftRegs_validOut_0 <= shiftRegs_validIn_delay_254_0;
      shiftRegs_validOut_1 <= shiftRegs_validIn_delay_254_1;
      shiftRegs_validOut_delay_1_0 <= shiftRegs_validOut_0;
      shiftRegs_validOut_delay_1_1 <= shiftRegs_validOut_1;
      shiftRegs_validOut_delay_2_0 <= shiftRegs_validOut_delay_1_0;
      shiftRegs_validOut_delay_2_1 <= shiftRegs_validOut_delay_1_1;
      shiftRegs_validOut_delay_3_0 <= shiftRegs_validOut_delay_2_0;
      shiftRegs_validOut_delay_3_1 <= shiftRegs_validOut_delay_2_1;
      shiftRegs_validOut_delay_4_0 <= shiftRegs_validOut_delay_3_0;
      shiftRegs_validOut_delay_4_1 <= shiftRegs_validOut_delay_3_1;
      shiftRegs_validOutFull_0 <= shiftRegs_validOut_delay_4_0;
      shiftRegs_validOutFull_1 <= shiftRegs_validOut_delay_4_1;
      if(io_dataOut_ready) begin
        outputValid <= 1'b0;
      end
      flushing_flushCnt_value <= flushing_flushCnt_valueNext;
      flushing_flushCnt_willOverflowIfInc <= (flushing_flushCnt_valueNext == 16'h9fff);
      stage1_NCnt_value <= stage1_NCnt_valueNext;
      stage1_NCnt_willOverflowIfInc <= (stage1_NCnt_valueNext == 32'hffffffff);
      stage1_GCnt_value <= stage1_GCnt_valueNext;
      stage1_GCnt_willOverflowIfInc <= (stage1_GCnt_valueNext == 4'b1001);
      stage1_emptyCnt_value <= stage1_emptyCnt_valueNext;
      stage1_emptyCnt_willOverflowIfInc <= (stage1_emptyCnt_valueNext == 9'h127);
      _zz_stage1_inputValid_0 <= (((((fsm_stateReg & fsm_enumDef_stage1) != 5'b00000) && (! stage1_waitReg)) && dataInBuffer_bufferOut_valid) && (_zz__zz_stage1_inputValid_0 != 13'h0));
      _zz_stage1_inputValid_0_1 <= _zz_stage1_inputValid_0;
      _zz_stage1_inputValid_0_2 <= _zz_stage1_inputValid_0_1;
      _zz_stage1_inputValid_0_3 <= _zz_stage1_inputValid_0_2;
      _zz_stage1_inputValid_0_4 <= _zz_stage1_inputValid_0_3;
      stage1_inputValid_0 <= _zz_stage1_inputValid_0_4;
      _zz_stage1_inputValid_1 <= (((((fsm_stateReg & fsm_enumDef_stage1) != 5'b00000) && (! stage1_waitReg)) && dataInBuffer_bufferOut_valid) && (_zz__zz_stage1_inputValid_1 != 13'h0));
      _zz_stage1_inputValid_1_1 <= _zz_stage1_inputValid_1;
      _zz_stage1_inputValid_1_2 <= _zz_stage1_inputValid_1_1;
      _zz_stage1_inputValid_1_3 <= _zz_stage1_inputValid_1_2;
      _zz_stage1_inputValid_1_4 <= _zz_stage1_inputValid_1_3;
      stage1_inputValid_1 <= _zz_stage1_inputValid_1_4;
      stage2_wCnt_value <= stage2_wCnt_valueNext;
      stage2_wCnt_willUnderflowIfDec <= (stage2_wCnt_valueNext == 12'h0);
      stage2_GCnt_value <= stage2_GCnt_valueNext;
      stage2_GCnt_willOverflowIfInc <= (stage2_GCnt_valueNext == 4'b1001);
      stage2_calCnt_value <= stage2_calCnt_valueNext;
      stage2_calCnt_willUnderflowIfDec <= (stage2_calCnt_valueNext == 2'b00);
      stage2_waitCnt_value <= stage2_waitCnt_valueNext;
      stage2_waitCnt_willOverflowIfInc <= (stage2_waitCnt_valueNext == 9'h125);
      stage3_GCnt_value <= stage3_GCnt_valueNext;
      stage3_GCnt_willUnderflowIfDec <= (stage3_GCnt_valueNext == 4'b0001);
      stage3_doubleCnt_value <= stage3_doubleCnt_valueNext;
      stage3_doubleCnt_willOverflowIfInc <= (stage3_doubleCnt_valueNext == 5'h19);
      stage3_doubleWaitCnt_value <= stage3_doubleWaitCnt_valueNext;
      stage3_doubleWaitCnt_willOverflowIfInc <= (stage3_doubleWaitCnt_valueNext == 9'h127);
      stage3_addWaitCnt_value <= stage3_addWaitCnt_valueNext;
      stage3_addWaitCnt_willOverflowIfInc <= (stage3_addWaitCnt_valueNext == 9'h127);
      stage3Final_doubleCnt_value <= stage3Final_doubleCnt_valueNext;
      stage3Final_doubleCnt_willOverflowIfInc <= (stage3Final_doubleCnt_valueNext == 4'b1100);
      stage3Final_doubleWaitCnt_value <= stage3Final_doubleWaitCnt_valueNext;
      stage3Final_doubleWaitCnt_willOverflowIfInc <= (stage3Final_doubleWaitCnt_valueNext == 9'h127);
      stage3Final_addWaitCnt_value <= stage3Final_addWaitCnt_valueNext;
      stage3Final_addWaitCnt_willOverflowIfInc <= (stage3Final_addWaitCnt_valueNext == 9'h127);
      fsm_stateReg <= fsm_stateNext;
      (* parallel_case *)
      case(1) // synthesis parallel_case
        (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
          if(when_Pippenger_l153) begin
            if(dataInBuffer_bufferOut_valid) begin
              if(stage1_GCnt_willOverflowIfInc) begin
                if(dataInBuffer_bufferOut_payload_last) begin
                  stage1_waitReg <= 1'b1;
                end
              end
              stage1_needAdd1_0 <= (|stage1_inputBarrelID_1[13 : 12]);
            end
          end else begin
            if(!when_Pippenger_l168) begin
              if(stage1_emptyCnt_willOverflowIfInc) begin
                stage1_waitReg <= 1'b0;
              end
            end
          end
        end
        (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
          if(when_Pippenger_l207) begin
            if(stage2_calCnt_willUnderflowIfDec) begin
              if(stage2_GCnt_willOverflowIfInc) begin
                stage2_waitReg <= 1'b1;
              end
            end
          end else begin
            if(stage2_waitCnt_willOverflowIfInc) begin
              stage2_waitReg <= 1'b0;
            end
          end
        end
        (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
          if(when_Pippenger_l249) begin
            if(stage3_doubleWaitCnt_willOverflowIfInc) begin
              if(stage3_doubleCnt_willOverflowIfInc) begin
                stage3_addReg <= 1'b1;
              end
            end
          end else begin
            if(stage3_addWaitCnt_willOverflowIfInc) begin
              stage3_addReg <= 1'b0;
            end
          end
        end
        (((fsm_stateReg) & fsm_enumDef_stage3Final) == fsm_enumDef_stage3Final) : begin
          if(when_Pippenger_l306) begin
            if(stage3Final_doubleWaitCnt_willOverflowIfInc) begin
              if(stage3Final_doubleCnt_willOverflowIfInc) begin
                stage3Final_addReg <= 1'b1;
              end
            end
          end else begin
            if(stage3Final_addWaitCnt_willOverflowIfInc) begin
              stage3Final_addReg <= 1'b0;
              stage3Final_pAddShr <= stage3Final_pAddShr[0 : 0];
              if(when_Pippenger_l319) begin
                outputValid <= 1'b1;
              end
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if(io_dataIn_ready) begin
      dataInBuffer_dataReg_last <= io_dataIn_payload_last;
      dataInBuffer_dataReg_fragment_P_X <= io_dataIn_payload_fragment_P_X;
      dataInBuffer_dataReg_fragment_P_Y <= io_dataIn_payload_fragment_P_Y;
      dataInBuffer_dataReg_fragment_P_Z <= io_dataIn_payload_fragment_P_Z;
      dataInBuffer_dataReg_fragment_P_T <= io_dataIn_payload_fragment_P_T;
      dataInBuffer_dataReg_fragment_K <= io_dataIn_payload_fragment_K;
    end else begin
      if(dataInBuffer_shift) begin
        dataInBuffer_dataReg_fragment_K <= {26'd0, _zz_dataInBuffer_dataReg_fragment_K};
      end
    end
    shiftRegs_addressIn_delay_1_0 <= shiftRegs_addressIn_0;
    shiftRegs_addressIn_delay_1_1 <= shiftRegs_addressIn_1;
    shiftRegs_addressIn_delay_2_0 <= shiftRegs_addressIn_delay_1_0;
    shiftRegs_addressIn_delay_2_1 <= shiftRegs_addressIn_delay_1_1;
    shiftRegs_addressIn_delay_3_0 <= shiftRegs_addressIn_delay_2_0;
    shiftRegs_addressIn_delay_3_1 <= shiftRegs_addressIn_delay_2_1;
    shiftRegs_addressIn_delay_4_0 <= shiftRegs_addressIn_delay_3_0;
    shiftRegs_addressIn_delay_4_1 <= shiftRegs_addressIn_delay_3_1;
    shiftRegs_addressIn_delay_5_0 <= shiftRegs_addressIn_delay_4_0;
    shiftRegs_addressIn_delay_5_1 <= shiftRegs_addressIn_delay_4_1;
    shiftRegs_addressIn_delay_6_0 <= shiftRegs_addressIn_delay_5_0;
    shiftRegs_addressIn_delay_6_1 <= shiftRegs_addressIn_delay_5_1;
    shiftRegs_addressIn_delay_7_0 <= shiftRegs_addressIn_delay_6_0;
    shiftRegs_addressIn_delay_7_1 <= shiftRegs_addressIn_delay_6_1;
    shiftRegs_addressIn_delay_8_0 <= shiftRegs_addressIn_delay_7_0;
    shiftRegs_addressIn_delay_8_1 <= shiftRegs_addressIn_delay_7_1;
    shiftRegs_addressIn_delay_9_0 <= shiftRegs_addressIn_delay_8_0;
    shiftRegs_addressIn_delay_9_1 <= shiftRegs_addressIn_delay_8_1;
    shiftRegs_addressIn_delay_10_0 <= shiftRegs_addressIn_delay_9_0;
    shiftRegs_addressIn_delay_10_1 <= shiftRegs_addressIn_delay_9_1;
    shiftRegs_addressIn_delay_11_0 <= shiftRegs_addressIn_delay_10_0;
    shiftRegs_addressIn_delay_11_1 <= shiftRegs_addressIn_delay_10_1;
    shiftRegs_addressIn_delay_12_0 <= shiftRegs_addressIn_delay_11_0;
    shiftRegs_addressIn_delay_12_1 <= shiftRegs_addressIn_delay_11_1;
    shiftRegs_addressIn_delay_13_0 <= shiftRegs_addressIn_delay_12_0;
    shiftRegs_addressIn_delay_13_1 <= shiftRegs_addressIn_delay_12_1;
    shiftRegs_addressIn_delay_14_0 <= shiftRegs_addressIn_delay_13_0;
    shiftRegs_addressIn_delay_14_1 <= shiftRegs_addressIn_delay_13_1;
    shiftRegs_addressIn_delay_15_0 <= shiftRegs_addressIn_delay_14_0;
    shiftRegs_addressIn_delay_15_1 <= shiftRegs_addressIn_delay_14_1;
    shiftRegs_addressIn_delay_16_0 <= shiftRegs_addressIn_delay_15_0;
    shiftRegs_addressIn_delay_16_1 <= shiftRegs_addressIn_delay_15_1;
    shiftRegs_addressIn_delay_17_0 <= shiftRegs_addressIn_delay_16_0;
    shiftRegs_addressIn_delay_17_1 <= shiftRegs_addressIn_delay_16_1;
    shiftRegs_addressIn_delay_18_0 <= shiftRegs_addressIn_delay_17_0;
    shiftRegs_addressIn_delay_18_1 <= shiftRegs_addressIn_delay_17_1;
    shiftRegs_addressIn_delay_19_0 <= shiftRegs_addressIn_delay_18_0;
    shiftRegs_addressIn_delay_19_1 <= shiftRegs_addressIn_delay_18_1;
    shiftRegs_addressIn_delay_20_0 <= shiftRegs_addressIn_delay_19_0;
    shiftRegs_addressIn_delay_20_1 <= shiftRegs_addressIn_delay_19_1;
    shiftRegs_addressIn_delay_21_0 <= shiftRegs_addressIn_delay_20_0;
    shiftRegs_addressIn_delay_21_1 <= shiftRegs_addressIn_delay_20_1;
    shiftRegs_addressIn_delay_22_0 <= shiftRegs_addressIn_delay_21_0;
    shiftRegs_addressIn_delay_22_1 <= shiftRegs_addressIn_delay_21_1;
    shiftRegs_addressIn_delay_23_0 <= shiftRegs_addressIn_delay_22_0;
    shiftRegs_addressIn_delay_23_1 <= shiftRegs_addressIn_delay_22_1;
    shiftRegs_addressIn_delay_24_0 <= shiftRegs_addressIn_delay_23_0;
    shiftRegs_addressIn_delay_24_1 <= shiftRegs_addressIn_delay_23_1;
    shiftRegs_addressIn_delay_25_0 <= shiftRegs_addressIn_delay_24_0;
    shiftRegs_addressIn_delay_25_1 <= shiftRegs_addressIn_delay_24_1;
    shiftRegs_addressIn_delay_26_0 <= shiftRegs_addressIn_delay_25_0;
    shiftRegs_addressIn_delay_26_1 <= shiftRegs_addressIn_delay_25_1;
    shiftRegs_addressIn_delay_27_0 <= shiftRegs_addressIn_delay_26_0;
    shiftRegs_addressIn_delay_27_1 <= shiftRegs_addressIn_delay_26_1;
    shiftRegs_addressIn_delay_28_0 <= shiftRegs_addressIn_delay_27_0;
    shiftRegs_addressIn_delay_28_1 <= shiftRegs_addressIn_delay_27_1;
    shiftRegs_addressIn_delay_29_0 <= shiftRegs_addressIn_delay_28_0;
    shiftRegs_addressIn_delay_29_1 <= shiftRegs_addressIn_delay_28_1;
    shiftRegs_addressIn_delay_30_0 <= shiftRegs_addressIn_delay_29_0;
    shiftRegs_addressIn_delay_30_1 <= shiftRegs_addressIn_delay_29_1;
    shiftRegs_addressIn_delay_31_0 <= shiftRegs_addressIn_delay_30_0;
    shiftRegs_addressIn_delay_31_1 <= shiftRegs_addressIn_delay_30_1;
    shiftRegs_addressIn_delay_32_0 <= shiftRegs_addressIn_delay_31_0;
    shiftRegs_addressIn_delay_32_1 <= shiftRegs_addressIn_delay_31_1;
    shiftRegs_addressIn_delay_33_0 <= shiftRegs_addressIn_delay_32_0;
    shiftRegs_addressIn_delay_33_1 <= shiftRegs_addressIn_delay_32_1;
    shiftRegs_addressIn_delay_34_0 <= shiftRegs_addressIn_delay_33_0;
    shiftRegs_addressIn_delay_34_1 <= shiftRegs_addressIn_delay_33_1;
    shiftRegs_addressIn_delay_35_0 <= shiftRegs_addressIn_delay_34_0;
    shiftRegs_addressIn_delay_35_1 <= shiftRegs_addressIn_delay_34_1;
    shiftRegs_addressIn_delay_36_0 <= shiftRegs_addressIn_delay_35_0;
    shiftRegs_addressIn_delay_36_1 <= shiftRegs_addressIn_delay_35_1;
    shiftRegs_addressIn_delay_37_0 <= shiftRegs_addressIn_delay_36_0;
    shiftRegs_addressIn_delay_37_1 <= shiftRegs_addressIn_delay_36_1;
    shiftRegs_addressIn_delay_38_0 <= shiftRegs_addressIn_delay_37_0;
    shiftRegs_addressIn_delay_38_1 <= shiftRegs_addressIn_delay_37_1;
    shiftRegs_addressIn_delay_39_0 <= shiftRegs_addressIn_delay_38_0;
    shiftRegs_addressIn_delay_39_1 <= shiftRegs_addressIn_delay_38_1;
    shiftRegs_addressIn_delay_40_0 <= shiftRegs_addressIn_delay_39_0;
    shiftRegs_addressIn_delay_40_1 <= shiftRegs_addressIn_delay_39_1;
    shiftRegs_addressIn_delay_41_0 <= shiftRegs_addressIn_delay_40_0;
    shiftRegs_addressIn_delay_41_1 <= shiftRegs_addressIn_delay_40_1;
    shiftRegs_addressIn_delay_42_0 <= shiftRegs_addressIn_delay_41_0;
    shiftRegs_addressIn_delay_42_1 <= shiftRegs_addressIn_delay_41_1;
    shiftRegs_addressIn_delay_43_0 <= shiftRegs_addressIn_delay_42_0;
    shiftRegs_addressIn_delay_43_1 <= shiftRegs_addressIn_delay_42_1;
    shiftRegs_addressIn_delay_44_0 <= shiftRegs_addressIn_delay_43_0;
    shiftRegs_addressIn_delay_44_1 <= shiftRegs_addressIn_delay_43_1;
    shiftRegs_addressIn_delay_45_0 <= shiftRegs_addressIn_delay_44_0;
    shiftRegs_addressIn_delay_45_1 <= shiftRegs_addressIn_delay_44_1;
    shiftRegs_addressIn_delay_46_0 <= shiftRegs_addressIn_delay_45_0;
    shiftRegs_addressIn_delay_46_1 <= shiftRegs_addressIn_delay_45_1;
    shiftRegs_addressIn_delay_47_0 <= shiftRegs_addressIn_delay_46_0;
    shiftRegs_addressIn_delay_47_1 <= shiftRegs_addressIn_delay_46_1;
    shiftRegs_addressIn_delay_48_0 <= shiftRegs_addressIn_delay_47_0;
    shiftRegs_addressIn_delay_48_1 <= shiftRegs_addressIn_delay_47_1;
    shiftRegs_addressIn_delay_49_0 <= shiftRegs_addressIn_delay_48_0;
    shiftRegs_addressIn_delay_49_1 <= shiftRegs_addressIn_delay_48_1;
    shiftRegs_addressIn_delay_50_0 <= shiftRegs_addressIn_delay_49_0;
    shiftRegs_addressIn_delay_50_1 <= shiftRegs_addressIn_delay_49_1;
    shiftRegs_addressIn_delay_51_0 <= shiftRegs_addressIn_delay_50_0;
    shiftRegs_addressIn_delay_51_1 <= shiftRegs_addressIn_delay_50_1;
    shiftRegs_addressIn_delay_52_0 <= shiftRegs_addressIn_delay_51_0;
    shiftRegs_addressIn_delay_52_1 <= shiftRegs_addressIn_delay_51_1;
    shiftRegs_addressIn_delay_53_0 <= shiftRegs_addressIn_delay_52_0;
    shiftRegs_addressIn_delay_53_1 <= shiftRegs_addressIn_delay_52_1;
    shiftRegs_addressIn_delay_54_0 <= shiftRegs_addressIn_delay_53_0;
    shiftRegs_addressIn_delay_54_1 <= shiftRegs_addressIn_delay_53_1;
    shiftRegs_addressIn_delay_55_0 <= shiftRegs_addressIn_delay_54_0;
    shiftRegs_addressIn_delay_55_1 <= shiftRegs_addressIn_delay_54_1;
    shiftRegs_addressIn_delay_56_0 <= shiftRegs_addressIn_delay_55_0;
    shiftRegs_addressIn_delay_56_1 <= shiftRegs_addressIn_delay_55_1;
    shiftRegs_addressIn_delay_57_0 <= shiftRegs_addressIn_delay_56_0;
    shiftRegs_addressIn_delay_57_1 <= shiftRegs_addressIn_delay_56_1;
    shiftRegs_addressIn_delay_58_0 <= shiftRegs_addressIn_delay_57_0;
    shiftRegs_addressIn_delay_58_1 <= shiftRegs_addressIn_delay_57_1;
    shiftRegs_addressIn_delay_59_0 <= shiftRegs_addressIn_delay_58_0;
    shiftRegs_addressIn_delay_59_1 <= shiftRegs_addressIn_delay_58_1;
    shiftRegs_addressIn_delay_60_0 <= shiftRegs_addressIn_delay_59_0;
    shiftRegs_addressIn_delay_60_1 <= shiftRegs_addressIn_delay_59_1;
    shiftRegs_addressIn_delay_61_0 <= shiftRegs_addressIn_delay_60_0;
    shiftRegs_addressIn_delay_61_1 <= shiftRegs_addressIn_delay_60_1;
    shiftRegs_addressIn_delay_62_0 <= shiftRegs_addressIn_delay_61_0;
    shiftRegs_addressIn_delay_62_1 <= shiftRegs_addressIn_delay_61_1;
    shiftRegs_addressIn_delay_63_0 <= shiftRegs_addressIn_delay_62_0;
    shiftRegs_addressIn_delay_63_1 <= shiftRegs_addressIn_delay_62_1;
    shiftRegs_addressIn_delay_64_0 <= shiftRegs_addressIn_delay_63_0;
    shiftRegs_addressIn_delay_64_1 <= shiftRegs_addressIn_delay_63_1;
    shiftRegs_addressIn_delay_65_0 <= shiftRegs_addressIn_delay_64_0;
    shiftRegs_addressIn_delay_65_1 <= shiftRegs_addressIn_delay_64_1;
    shiftRegs_addressIn_delay_66_0 <= shiftRegs_addressIn_delay_65_0;
    shiftRegs_addressIn_delay_66_1 <= shiftRegs_addressIn_delay_65_1;
    shiftRegs_addressIn_delay_67_0 <= shiftRegs_addressIn_delay_66_0;
    shiftRegs_addressIn_delay_67_1 <= shiftRegs_addressIn_delay_66_1;
    shiftRegs_addressIn_delay_68_0 <= shiftRegs_addressIn_delay_67_0;
    shiftRegs_addressIn_delay_68_1 <= shiftRegs_addressIn_delay_67_1;
    shiftRegs_addressIn_delay_69_0 <= shiftRegs_addressIn_delay_68_0;
    shiftRegs_addressIn_delay_69_1 <= shiftRegs_addressIn_delay_68_1;
    shiftRegs_addressIn_delay_70_0 <= shiftRegs_addressIn_delay_69_0;
    shiftRegs_addressIn_delay_70_1 <= shiftRegs_addressIn_delay_69_1;
    shiftRegs_addressIn_delay_71_0 <= shiftRegs_addressIn_delay_70_0;
    shiftRegs_addressIn_delay_71_1 <= shiftRegs_addressIn_delay_70_1;
    shiftRegs_addressIn_delay_72_0 <= shiftRegs_addressIn_delay_71_0;
    shiftRegs_addressIn_delay_72_1 <= shiftRegs_addressIn_delay_71_1;
    shiftRegs_addressIn_delay_73_0 <= shiftRegs_addressIn_delay_72_0;
    shiftRegs_addressIn_delay_73_1 <= shiftRegs_addressIn_delay_72_1;
    shiftRegs_addressIn_delay_74_0 <= shiftRegs_addressIn_delay_73_0;
    shiftRegs_addressIn_delay_74_1 <= shiftRegs_addressIn_delay_73_1;
    shiftRegs_addressIn_delay_75_0 <= shiftRegs_addressIn_delay_74_0;
    shiftRegs_addressIn_delay_75_1 <= shiftRegs_addressIn_delay_74_1;
    shiftRegs_addressIn_delay_76_0 <= shiftRegs_addressIn_delay_75_0;
    shiftRegs_addressIn_delay_76_1 <= shiftRegs_addressIn_delay_75_1;
    shiftRegs_addressIn_delay_77_0 <= shiftRegs_addressIn_delay_76_0;
    shiftRegs_addressIn_delay_77_1 <= shiftRegs_addressIn_delay_76_1;
    shiftRegs_addressIn_delay_78_0 <= shiftRegs_addressIn_delay_77_0;
    shiftRegs_addressIn_delay_78_1 <= shiftRegs_addressIn_delay_77_1;
    shiftRegs_addressIn_delay_79_0 <= shiftRegs_addressIn_delay_78_0;
    shiftRegs_addressIn_delay_79_1 <= shiftRegs_addressIn_delay_78_1;
    shiftRegs_addressIn_delay_80_0 <= shiftRegs_addressIn_delay_79_0;
    shiftRegs_addressIn_delay_80_1 <= shiftRegs_addressIn_delay_79_1;
    shiftRegs_addressIn_delay_81_0 <= shiftRegs_addressIn_delay_80_0;
    shiftRegs_addressIn_delay_81_1 <= shiftRegs_addressIn_delay_80_1;
    shiftRegs_addressIn_delay_82_0 <= shiftRegs_addressIn_delay_81_0;
    shiftRegs_addressIn_delay_82_1 <= shiftRegs_addressIn_delay_81_1;
    shiftRegs_addressIn_delay_83_0 <= shiftRegs_addressIn_delay_82_0;
    shiftRegs_addressIn_delay_83_1 <= shiftRegs_addressIn_delay_82_1;
    shiftRegs_addressIn_delay_84_0 <= shiftRegs_addressIn_delay_83_0;
    shiftRegs_addressIn_delay_84_1 <= shiftRegs_addressIn_delay_83_1;
    shiftRegs_addressIn_delay_85_0 <= shiftRegs_addressIn_delay_84_0;
    shiftRegs_addressIn_delay_85_1 <= shiftRegs_addressIn_delay_84_1;
    shiftRegs_addressIn_delay_86_0 <= shiftRegs_addressIn_delay_85_0;
    shiftRegs_addressIn_delay_86_1 <= shiftRegs_addressIn_delay_85_1;
    shiftRegs_addressIn_delay_87_0 <= shiftRegs_addressIn_delay_86_0;
    shiftRegs_addressIn_delay_87_1 <= shiftRegs_addressIn_delay_86_1;
    shiftRegs_addressIn_delay_88_0 <= shiftRegs_addressIn_delay_87_0;
    shiftRegs_addressIn_delay_88_1 <= shiftRegs_addressIn_delay_87_1;
    shiftRegs_addressIn_delay_89_0 <= shiftRegs_addressIn_delay_88_0;
    shiftRegs_addressIn_delay_89_1 <= shiftRegs_addressIn_delay_88_1;
    shiftRegs_addressIn_delay_90_0 <= shiftRegs_addressIn_delay_89_0;
    shiftRegs_addressIn_delay_90_1 <= shiftRegs_addressIn_delay_89_1;
    shiftRegs_addressIn_delay_91_0 <= shiftRegs_addressIn_delay_90_0;
    shiftRegs_addressIn_delay_91_1 <= shiftRegs_addressIn_delay_90_1;
    shiftRegs_addressIn_delay_92_0 <= shiftRegs_addressIn_delay_91_0;
    shiftRegs_addressIn_delay_92_1 <= shiftRegs_addressIn_delay_91_1;
    shiftRegs_addressIn_delay_93_0 <= shiftRegs_addressIn_delay_92_0;
    shiftRegs_addressIn_delay_93_1 <= shiftRegs_addressIn_delay_92_1;
    shiftRegs_addressIn_delay_94_0 <= shiftRegs_addressIn_delay_93_0;
    shiftRegs_addressIn_delay_94_1 <= shiftRegs_addressIn_delay_93_1;
    shiftRegs_addressIn_delay_95_0 <= shiftRegs_addressIn_delay_94_0;
    shiftRegs_addressIn_delay_95_1 <= shiftRegs_addressIn_delay_94_1;
    shiftRegs_addressIn_delay_96_0 <= shiftRegs_addressIn_delay_95_0;
    shiftRegs_addressIn_delay_96_1 <= shiftRegs_addressIn_delay_95_1;
    shiftRegs_addressIn_delay_97_0 <= shiftRegs_addressIn_delay_96_0;
    shiftRegs_addressIn_delay_97_1 <= shiftRegs_addressIn_delay_96_1;
    shiftRegs_addressIn_delay_98_0 <= shiftRegs_addressIn_delay_97_0;
    shiftRegs_addressIn_delay_98_1 <= shiftRegs_addressIn_delay_97_1;
    shiftRegs_addressIn_delay_99_0 <= shiftRegs_addressIn_delay_98_0;
    shiftRegs_addressIn_delay_99_1 <= shiftRegs_addressIn_delay_98_1;
    shiftRegs_addressIn_delay_100_0 <= shiftRegs_addressIn_delay_99_0;
    shiftRegs_addressIn_delay_100_1 <= shiftRegs_addressIn_delay_99_1;
    shiftRegs_addressIn_delay_101_0 <= shiftRegs_addressIn_delay_100_0;
    shiftRegs_addressIn_delay_101_1 <= shiftRegs_addressIn_delay_100_1;
    shiftRegs_addressIn_delay_102_0 <= shiftRegs_addressIn_delay_101_0;
    shiftRegs_addressIn_delay_102_1 <= shiftRegs_addressIn_delay_101_1;
    shiftRegs_addressIn_delay_103_0 <= shiftRegs_addressIn_delay_102_0;
    shiftRegs_addressIn_delay_103_1 <= shiftRegs_addressIn_delay_102_1;
    shiftRegs_addressIn_delay_104_0 <= shiftRegs_addressIn_delay_103_0;
    shiftRegs_addressIn_delay_104_1 <= shiftRegs_addressIn_delay_103_1;
    shiftRegs_addressIn_delay_105_0 <= shiftRegs_addressIn_delay_104_0;
    shiftRegs_addressIn_delay_105_1 <= shiftRegs_addressIn_delay_104_1;
    shiftRegs_addressIn_delay_106_0 <= shiftRegs_addressIn_delay_105_0;
    shiftRegs_addressIn_delay_106_1 <= shiftRegs_addressIn_delay_105_1;
    shiftRegs_addressIn_delay_107_0 <= shiftRegs_addressIn_delay_106_0;
    shiftRegs_addressIn_delay_107_1 <= shiftRegs_addressIn_delay_106_1;
    shiftRegs_addressIn_delay_108_0 <= shiftRegs_addressIn_delay_107_0;
    shiftRegs_addressIn_delay_108_1 <= shiftRegs_addressIn_delay_107_1;
    shiftRegs_addressIn_delay_109_0 <= shiftRegs_addressIn_delay_108_0;
    shiftRegs_addressIn_delay_109_1 <= shiftRegs_addressIn_delay_108_1;
    shiftRegs_addressIn_delay_110_0 <= shiftRegs_addressIn_delay_109_0;
    shiftRegs_addressIn_delay_110_1 <= shiftRegs_addressIn_delay_109_1;
    shiftRegs_addressIn_delay_111_0 <= shiftRegs_addressIn_delay_110_0;
    shiftRegs_addressIn_delay_111_1 <= shiftRegs_addressIn_delay_110_1;
    shiftRegs_addressIn_delay_112_0 <= shiftRegs_addressIn_delay_111_0;
    shiftRegs_addressIn_delay_112_1 <= shiftRegs_addressIn_delay_111_1;
    shiftRegs_addressIn_delay_113_0 <= shiftRegs_addressIn_delay_112_0;
    shiftRegs_addressIn_delay_113_1 <= shiftRegs_addressIn_delay_112_1;
    shiftRegs_addressIn_delay_114_0 <= shiftRegs_addressIn_delay_113_0;
    shiftRegs_addressIn_delay_114_1 <= shiftRegs_addressIn_delay_113_1;
    shiftRegs_addressIn_delay_115_0 <= shiftRegs_addressIn_delay_114_0;
    shiftRegs_addressIn_delay_115_1 <= shiftRegs_addressIn_delay_114_1;
    shiftRegs_addressIn_delay_116_0 <= shiftRegs_addressIn_delay_115_0;
    shiftRegs_addressIn_delay_116_1 <= shiftRegs_addressIn_delay_115_1;
    shiftRegs_addressIn_delay_117_0 <= shiftRegs_addressIn_delay_116_0;
    shiftRegs_addressIn_delay_117_1 <= shiftRegs_addressIn_delay_116_1;
    shiftRegs_addressIn_delay_118_0 <= shiftRegs_addressIn_delay_117_0;
    shiftRegs_addressIn_delay_118_1 <= shiftRegs_addressIn_delay_117_1;
    shiftRegs_addressIn_delay_119_0 <= shiftRegs_addressIn_delay_118_0;
    shiftRegs_addressIn_delay_119_1 <= shiftRegs_addressIn_delay_118_1;
    shiftRegs_addressIn_delay_120_0 <= shiftRegs_addressIn_delay_119_0;
    shiftRegs_addressIn_delay_120_1 <= shiftRegs_addressIn_delay_119_1;
    shiftRegs_addressIn_delay_121_0 <= shiftRegs_addressIn_delay_120_0;
    shiftRegs_addressIn_delay_121_1 <= shiftRegs_addressIn_delay_120_1;
    shiftRegs_addressIn_delay_122_0 <= shiftRegs_addressIn_delay_121_0;
    shiftRegs_addressIn_delay_122_1 <= shiftRegs_addressIn_delay_121_1;
    shiftRegs_addressIn_delay_123_0 <= shiftRegs_addressIn_delay_122_0;
    shiftRegs_addressIn_delay_123_1 <= shiftRegs_addressIn_delay_122_1;
    shiftRegs_addressIn_delay_124_0 <= shiftRegs_addressIn_delay_123_0;
    shiftRegs_addressIn_delay_124_1 <= shiftRegs_addressIn_delay_123_1;
    shiftRegs_addressIn_delay_125_0 <= shiftRegs_addressIn_delay_124_0;
    shiftRegs_addressIn_delay_125_1 <= shiftRegs_addressIn_delay_124_1;
    shiftRegs_addressIn_delay_126_0 <= shiftRegs_addressIn_delay_125_0;
    shiftRegs_addressIn_delay_126_1 <= shiftRegs_addressIn_delay_125_1;
    shiftRegs_addressIn_delay_127_0 <= shiftRegs_addressIn_delay_126_0;
    shiftRegs_addressIn_delay_127_1 <= shiftRegs_addressIn_delay_126_1;
    shiftRegs_addressIn_delay_128_0 <= shiftRegs_addressIn_delay_127_0;
    shiftRegs_addressIn_delay_128_1 <= shiftRegs_addressIn_delay_127_1;
    shiftRegs_addressIn_delay_129_0 <= shiftRegs_addressIn_delay_128_0;
    shiftRegs_addressIn_delay_129_1 <= shiftRegs_addressIn_delay_128_1;
    shiftRegs_addressIn_delay_130_0 <= shiftRegs_addressIn_delay_129_0;
    shiftRegs_addressIn_delay_130_1 <= shiftRegs_addressIn_delay_129_1;
    shiftRegs_addressIn_delay_131_0 <= shiftRegs_addressIn_delay_130_0;
    shiftRegs_addressIn_delay_131_1 <= shiftRegs_addressIn_delay_130_1;
    shiftRegs_addressIn_delay_132_0 <= shiftRegs_addressIn_delay_131_0;
    shiftRegs_addressIn_delay_132_1 <= shiftRegs_addressIn_delay_131_1;
    shiftRegs_addressIn_delay_133_0 <= shiftRegs_addressIn_delay_132_0;
    shiftRegs_addressIn_delay_133_1 <= shiftRegs_addressIn_delay_132_1;
    shiftRegs_addressIn_delay_134_0 <= shiftRegs_addressIn_delay_133_0;
    shiftRegs_addressIn_delay_134_1 <= shiftRegs_addressIn_delay_133_1;
    shiftRegs_addressIn_delay_135_0 <= shiftRegs_addressIn_delay_134_0;
    shiftRegs_addressIn_delay_135_1 <= shiftRegs_addressIn_delay_134_1;
    shiftRegs_addressIn_delay_136_0 <= shiftRegs_addressIn_delay_135_0;
    shiftRegs_addressIn_delay_136_1 <= shiftRegs_addressIn_delay_135_1;
    shiftRegs_addressIn_delay_137_0 <= shiftRegs_addressIn_delay_136_0;
    shiftRegs_addressIn_delay_137_1 <= shiftRegs_addressIn_delay_136_1;
    shiftRegs_addressIn_delay_138_0 <= shiftRegs_addressIn_delay_137_0;
    shiftRegs_addressIn_delay_138_1 <= shiftRegs_addressIn_delay_137_1;
    shiftRegs_addressIn_delay_139_0 <= shiftRegs_addressIn_delay_138_0;
    shiftRegs_addressIn_delay_139_1 <= shiftRegs_addressIn_delay_138_1;
    shiftRegs_addressIn_delay_140_0 <= shiftRegs_addressIn_delay_139_0;
    shiftRegs_addressIn_delay_140_1 <= shiftRegs_addressIn_delay_139_1;
    shiftRegs_addressIn_delay_141_0 <= shiftRegs_addressIn_delay_140_0;
    shiftRegs_addressIn_delay_141_1 <= shiftRegs_addressIn_delay_140_1;
    shiftRegs_addressIn_delay_142_0 <= shiftRegs_addressIn_delay_141_0;
    shiftRegs_addressIn_delay_142_1 <= shiftRegs_addressIn_delay_141_1;
    shiftRegs_addressIn_delay_143_0 <= shiftRegs_addressIn_delay_142_0;
    shiftRegs_addressIn_delay_143_1 <= shiftRegs_addressIn_delay_142_1;
    shiftRegs_addressIn_delay_144_0 <= shiftRegs_addressIn_delay_143_0;
    shiftRegs_addressIn_delay_144_1 <= shiftRegs_addressIn_delay_143_1;
    shiftRegs_addressIn_delay_145_0 <= shiftRegs_addressIn_delay_144_0;
    shiftRegs_addressIn_delay_145_1 <= shiftRegs_addressIn_delay_144_1;
    shiftRegs_addressIn_delay_146_0 <= shiftRegs_addressIn_delay_145_0;
    shiftRegs_addressIn_delay_146_1 <= shiftRegs_addressIn_delay_145_1;
    shiftRegs_addressIn_delay_147_0 <= shiftRegs_addressIn_delay_146_0;
    shiftRegs_addressIn_delay_147_1 <= shiftRegs_addressIn_delay_146_1;
    shiftRegs_addressIn_delay_148_0 <= shiftRegs_addressIn_delay_147_0;
    shiftRegs_addressIn_delay_148_1 <= shiftRegs_addressIn_delay_147_1;
    shiftRegs_addressIn_delay_149_0 <= shiftRegs_addressIn_delay_148_0;
    shiftRegs_addressIn_delay_149_1 <= shiftRegs_addressIn_delay_148_1;
    shiftRegs_addressIn_delay_150_0 <= shiftRegs_addressIn_delay_149_0;
    shiftRegs_addressIn_delay_150_1 <= shiftRegs_addressIn_delay_149_1;
    shiftRegs_addressIn_delay_151_0 <= shiftRegs_addressIn_delay_150_0;
    shiftRegs_addressIn_delay_151_1 <= shiftRegs_addressIn_delay_150_1;
    shiftRegs_addressIn_delay_152_0 <= shiftRegs_addressIn_delay_151_0;
    shiftRegs_addressIn_delay_152_1 <= shiftRegs_addressIn_delay_151_1;
    shiftRegs_addressIn_delay_153_0 <= shiftRegs_addressIn_delay_152_0;
    shiftRegs_addressIn_delay_153_1 <= shiftRegs_addressIn_delay_152_1;
    shiftRegs_addressIn_delay_154_0 <= shiftRegs_addressIn_delay_153_0;
    shiftRegs_addressIn_delay_154_1 <= shiftRegs_addressIn_delay_153_1;
    shiftRegs_addressIn_delay_155_0 <= shiftRegs_addressIn_delay_154_0;
    shiftRegs_addressIn_delay_155_1 <= shiftRegs_addressIn_delay_154_1;
    shiftRegs_addressIn_delay_156_0 <= shiftRegs_addressIn_delay_155_0;
    shiftRegs_addressIn_delay_156_1 <= shiftRegs_addressIn_delay_155_1;
    shiftRegs_addressIn_delay_157_0 <= shiftRegs_addressIn_delay_156_0;
    shiftRegs_addressIn_delay_157_1 <= shiftRegs_addressIn_delay_156_1;
    shiftRegs_addressIn_delay_158_0 <= shiftRegs_addressIn_delay_157_0;
    shiftRegs_addressIn_delay_158_1 <= shiftRegs_addressIn_delay_157_1;
    shiftRegs_addressIn_delay_159_0 <= shiftRegs_addressIn_delay_158_0;
    shiftRegs_addressIn_delay_159_1 <= shiftRegs_addressIn_delay_158_1;
    shiftRegs_addressIn_delay_160_0 <= shiftRegs_addressIn_delay_159_0;
    shiftRegs_addressIn_delay_160_1 <= shiftRegs_addressIn_delay_159_1;
    shiftRegs_addressIn_delay_161_0 <= shiftRegs_addressIn_delay_160_0;
    shiftRegs_addressIn_delay_161_1 <= shiftRegs_addressIn_delay_160_1;
    shiftRegs_addressIn_delay_162_0 <= shiftRegs_addressIn_delay_161_0;
    shiftRegs_addressIn_delay_162_1 <= shiftRegs_addressIn_delay_161_1;
    shiftRegs_addressIn_delay_163_0 <= shiftRegs_addressIn_delay_162_0;
    shiftRegs_addressIn_delay_163_1 <= shiftRegs_addressIn_delay_162_1;
    shiftRegs_addressIn_delay_164_0 <= shiftRegs_addressIn_delay_163_0;
    shiftRegs_addressIn_delay_164_1 <= shiftRegs_addressIn_delay_163_1;
    shiftRegs_addressIn_delay_165_0 <= shiftRegs_addressIn_delay_164_0;
    shiftRegs_addressIn_delay_165_1 <= shiftRegs_addressIn_delay_164_1;
    shiftRegs_addressIn_delay_166_0 <= shiftRegs_addressIn_delay_165_0;
    shiftRegs_addressIn_delay_166_1 <= shiftRegs_addressIn_delay_165_1;
    shiftRegs_addressIn_delay_167_0 <= shiftRegs_addressIn_delay_166_0;
    shiftRegs_addressIn_delay_167_1 <= shiftRegs_addressIn_delay_166_1;
    shiftRegs_addressIn_delay_168_0 <= shiftRegs_addressIn_delay_167_0;
    shiftRegs_addressIn_delay_168_1 <= shiftRegs_addressIn_delay_167_1;
    shiftRegs_addressIn_delay_169_0 <= shiftRegs_addressIn_delay_168_0;
    shiftRegs_addressIn_delay_169_1 <= shiftRegs_addressIn_delay_168_1;
    shiftRegs_addressIn_delay_170_0 <= shiftRegs_addressIn_delay_169_0;
    shiftRegs_addressIn_delay_170_1 <= shiftRegs_addressIn_delay_169_1;
    shiftRegs_addressIn_delay_171_0 <= shiftRegs_addressIn_delay_170_0;
    shiftRegs_addressIn_delay_171_1 <= shiftRegs_addressIn_delay_170_1;
    shiftRegs_addressIn_delay_172_0 <= shiftRegs_addressIn_delay_171_0;
    shiftRegs_addressIn_delay_172_1 <= shiftRegs_addressIn_delay_171_1;
    shiftRegs_addressIn_delay_173_0 <= shiftRegs_addressIn_delay_172_0;
    shiftRegs_addressIn_delay_173_1 <= shiftRegs_addressIn_delay_172_1;
    shiftRegs_addressIn_delay_174_0 <= shiftRegs_addressIn_delay_173_0;
    shiftRegs_addressIn_delay_174_1 <= shiftRegs_addressIn_delay_173_1;
    shiftRegs_addressIn_delay_175_0 <= shiftRegs_addressIn_delay_174_0;
    shiftRegs_addressIn_delay_175_1 <= shiftRegs_addressIn_delay_174_1;
    shiftRegs_addressIn_delay_176_0 <= shiftRegs_addressIn_delay_175_0;
    shiftRegs_addressIn_delay_176_1 <= shiftRegs_addressIn_delay_175_1;
    shiftRegs_addressIn_delay_177_0 <= shiftRegs_addressIn_delay_176_0;
    shiftRegs_addressIn_delay_177_1 <= shiftRegs_addressIn_delay_176_1;
    shiftRegs_addressIn_delay_178_0 <= shiftRegs_addressIn_delay_177_0;
    shiftRegs_addressIn_delay_178_1 <= shiftRegs_addressIn_delay_177_1;
    shiftRegs_addressIn_delay_179_0 <= shiftRegs_addressIn_delay_178_0;
    shiftRegs_addressIn_delay_179_1 <= shiftRegs_addressIn_delay_178_1;
    shiftRegs_addressIn_delay_180_0 <= shiftRegs_addressIn_delay_179_0;
    shiftRegs_addressIn_delay_180_1 <= shiftRegs_addressIn_delay_179_1;
    shiftRegs_addressIn_delay_181_0 <= shiftRegs_addressIn_delay_180_0;
    shiftRegs_addressIn_delay_181_1 <= shiftRegs_addressIn_delay_180_1;
    shiftRegs_addressIn_delay_182_0 <= shiftRegs_addressIn_delay_181_0;
    shiftRegs_addressIn_delay_182_1 <= shiftRegs_addressIn_delay_181_1;
    shiftRegs_addressIn_delay_183_0 <= shiftRegs_addressIn_delay_182_0;
    shiftRegs_addressIn_delay_183_1 <= shiftRegs_addressIn_delay_182_1;
    shiftRegs_addressIn_delay_184_0 <= shiftRegs_addressIn_delay_183_0;
    shiftRegs_addressIn_delay_184_1 <= shiftRegs_addressIn_delay_183_1;
    shiftRegs_addressIn_delay_185_0 <= shiftRegs_addressIn_delay_184_0;
    shiftRegs_addressIn_delay_185_1 <= shiftRegs_addressIn_delay_184_1;
    shiftRegs_addressIn_delay_186_0 <= shiftRegs_addressIn_delay_185_0;
    shiftRegs_addressIn_delay_186_1 <= shiftRegs_addressIn_delay_185_1;
    shiftRegs_addressIn_delay_187_0 <= shiftRegs_addressIn_delay_186_0;
    shiftRegs_addressIn_delay_187_1 <= shiftRegs_addressIn_delay_186_1;
    shiftRegs_addressIn_delay_188_0 <= shiftRegs_addressIn_delay_187_0;
    shiftRegs_addressIn_delay_188_1 <= shiftRegs_addressIn_delay_187_1;
    shiftRegs_addressIn_delay_189_0 <= shiftRegs_addressIn_delay_188_0;
    shiftRegs_addressIn_delay_189_1 <= shiftRegs_addressIn_delay_188_1;
    shiftRegs_addressIn_delay_190_0 <= shiftRegs_addressIn_delay_189_0;
    shiftRegs_addressIn_delay_190_1 <= shiftRegs_addressIn_delay_189_1;
    shiftRegs_addressIn_delay_191_0 <= shiftRegs_addressIn_delay_190_0;
    shiftRegs_addressIn_delay_191_1 <= shiftRegs_addressIn_delay_190_1;
    shiftRegs_addressIn_delay_192_0 <= shiftRegs_addressIn_delay_191_0;
    shiftRegs_addressIn_delay_192_1 <= shiftRegs_addressIn_delay_191_1;
    shiftRegs_addressIn_delay_193_0 <= shiftRegs_addressIn_delay_192_0;
    shiftRegs_addressIn_delay_193_1 <= shiftRegs_addressIn_delay_192_1;
    shiftRegs_addressIn_delay_194_0 <= shiftRegs_addressIn_delay_193_0;
    shiftRegs_addressIn_delay_194_1 <= shiftRegs_addressIn_delay_193_1;
    shiftRegs_addressIn_delay_195_0 <= shiftRegs_addressIn_delay_194_0;
    shiftRegs_addressIn_delay_195_1 <= shiftRegs_addressIn_delay_194_1;
    shiftRegs_addressIn_delay_196_0 <= shiftRegs_addressIn_delay_195_0;
    shiftRegs_addressIn_delay_196_1 <= shiftRegs_addressIn_delay_195_1;
    shiftRegs_addressIn_delay_197_0 <= shiftRegs_addressIn_delay_196_0;
    shiftRegs_addressIn_delay_197_1 <= shiftRegs_addressIn_delay_196_1;
    shiftRegs_addressIn_delay_198_0 <= shiftRegs_addressIn_delay_197_0;
    shiftRegs_addressIn_delay_198_1 <= shiftRegs_addressIn_delay_197_1;
    shiftRegs_addressIn_delay_199_0 <= shiftRegs_addressIn_delay_198_0;
    shiftRegs_addressIn_delay_199_1 <= shiftRegs_addressIn_delay_198_1;
    shiftRegs_addressIn_delay_200_0 <= shiftRegs_addressIn_delay_199_0;
    shiftRegs_addressIn_delay_200_1 <= shiftRegs_addressIn_delay_199_1;
    shiftRegs_addressIn_delay_201_0 <= shiftRegs_addressIn_delay_200_0;
    shiftRegs_addressIn_delay_201_1 <= shiftRegs_addressIn_delay_200_1;
    shiftRegs_addressIn_delay_202_0 <= shiftRegs_addressIn_delay_201_0;
    shiftRegs_addressIn_delay_202_1 <= shiftRegs_addressIn_delay_201_1;
    shiftRegs_addressIn_delay_203_0 <= shiftRegs_addressIn_delay_202_0;
    shiftRegs_addressIn_delay_203_1 <= shiftRegs_addressIn_delay_202_1;
    shiftRegs_addressIn_delay_204_0 <= shiftRegs_addressIn_delay_203_0;
    shiftRegs_addressIn_delay_204_1 <= shiftRegs_addressIn_delay_203_1;
    shiftRegs_addressIn_delay_205_0 <= shiftRegs_addressIn_delay_204_0;
    shiftRegs_addressIn_delay_205_1 <= shiftRegs_addressIn_delay_204_1;
    shiftRegs_addressIn_delay_206_0 <= shiftRegs_addressIn_delay_205_0;
    shiftRegs_addressIn_delay_206_1 <= shiftRegs_addressIn_delay_205_1;
    shiftRegs_addressIn_delay_207_0 <= shiftRegs_addressIn_delay_206_0;
    shiftRegs_addressIn_delay_207_1 <= shiftRegs_addressIn_delay_206_1;
    shiftRegs_addressIn_delay_208_0 <= shiftRegs_addressIn_delay_207_0;
    shiftRegs_addressIn_delay_208_1 <= shiftRegs_addressIn_delay_207_1;
    shiftRegs_addressIn_delay_209_0 <= shiftRegs_addressIn_delay_208_0;
    shiftRegs_addressIn_delay_209_1 <= shiftRegs_addressIn_delay_208_1;
    shiftRegs_addressIn_delay_210_0 <= shiftRegs_addressIn_delay_209_0;
    shiftRegs_addressIn_delay_210_1 <= shiftRegs_addressIn_delay_209_1;
    shiftRegs_addressIn_delay_211_0 <= shiftRegs_addressIn_delay_210_0;
    shiftRegs_addressIn_delay_211_1 <= shiftRegs_addressIn_delay_210_1;
    shiftRegs_addressIn_delay_212_0 <= shiftRegs_addressIn_delay_211_0;
    shiftRegs_addressIn_delay_212_1 <= shiftRegs_addressIn_delay_211_1;
    shiftRegs_addressIn_delay_213_0 <= shiftRegs_addressIn_delay_212_0;
    shiftRegs_addressIn_delay_213_1 <= shiftRegs_addressIn_delay_212_1;
    shiftRegs_addressIn_delay_214_0 <= shiftRegs_addressIn_delay_213_0;
    shiftRegs_addressIn_delay_214_1 <= shiftRegs_addressIn_delay_213_1;
    shiftRegs_addressIn_delay_215_0 <= shiftRegs_addressIn_delay_214_0;
    shiftRegs_addressIn_delay_215_1 <= shiftRegs_addressIn_delay_214_1;
    shiftRegs_addressIn_delay_216_0 <= shiftRegs_addressIn_delay_215_0;
    shiftRegs_addressIn_delay_216_1 <= shiftRegs_addressIn_delay_215_1;
    shiftRegs_addressIn_delay_217_0 <= shiftRegs_addressIn_delay_216_0;
    shiftRegs_addressIn_delay_217_1 <= shiftRegs_addressIn_delay_216_1;
    shiftRegs_addressIn_delay_218_0 <= shiftRegs_addressIn_delay_217_0;
    shiftRegs_addressIn_delay_218_1 <= shiftRegs_addressIn_delay_217_1;
    shiftRegs_addressIn_delay_219_0 <= shiftRegs_addressIn_delay_218_0;
    shiftRegs_addressIn_delay_219_1 <= shiftRegs_addressIn_delay_218_1;
    shiftRegs_addressIn_delay_220_0 <= shiftRegs_addressIn_delay_219_0;
    shiftRegs_addressIn_delay_220_1 <= shiftRegs_addressIn_delay_219_1;
    shiftRegs_addressIn_delay_221_0 <= shiftRegs_addressIn_delay_220_0;
    shiftRegs_addressIn_delay_221_1 <= shiftRegs_addressIn_delay_220_1;
    shiftRegs_addressIn_delay_222_0 <= shiftRegs_addressIn_delay_221_0;
    shiftRegs_addressIn_delay_222_1 <= shiftRegs_addressIn_delay_221_1;
    shiftRegs_addressIn_delay_223_0 <= shiftRegs_addressIn_delay_222_0;
    shiftRegs_addressIn_delay_223_1 <= shiftRegs_addressIn_delay_222_1;
    shiftRegs_addressIn_delay_224_0 <= shiftRegs_addressIn_delay_223_0;
    shiftRegs_addressIn_delay_224_1 <= shiftRegs_addressIn_delay_223_1;
    shiftRegs_addressIn_delay_225_0 <= shiftRegs_addressIn_delay_224_0;
    shiftRegs_addressIn_delay_225_1 <= shiftRegs_addressIn_delay_224_1;
    shiftRegs_addressIn_delay_226_0 <= shiftRegs_addressIn_delay_225_0;
    shiftRegs_addressIn_delay_226_1 <= shiftRegs_addressIn_delay_225_1;
    shiftRegs_addressIn_delay_227_0 <= shiftRegs_addressIn_delay_226_0;
    shiftRegs_addressIn_delay_227_1 <= shiftRegs_addressIn_delay_226_1;
    shiftRegs_addressIn_delay_228_0 <= shiftRegs_addressIn_delay_227_0;
    shiftRegs_addressIn_delay_228_1 <= shiftRegs_addressIn_delay_227_1;
    shiftRegs_addressIn_delay_229_0 <= shiftRegs_addressIn_delay_228_0;
    shiftRegs_addressIn_delay_229_1 <= shiftRegs_addressIn_delay_228_1;
    shiftRegs_addressIn_delay_230_0 <= shiftRegs_addressIn_delay_229_0;
    shiftRegs_addressIn_delay_230_1 <= shiftRegs_addressIn_delay_229_1;
    shiftRegs_addressIn_delay_231_0 <= shiftRegs_addressIn_delay_230_0;
    shiftRegs_addressIn_delay_231_1 <= shiftRegs_addressIn_delay_230_1;
    shiftRegs_addressIn_delay_232_0 <= shiftRegs_addressIn_delay_231_0;
    shiftRegs_addressIn_delay_232_1 <= shiftRegs_addressIn_delay_231_1;
    shiftRegs_addressIn_delay_233_0 <= shiftRegs_addressIn_delay_232_0;
    shiftRegs_addressIn_delay_233_1 <= shiftRegs_addressIn_delay_232_1;
    shiftRegs_addressIn_delay_234_0 <= shiftRegs_addressIn_delay_233_0;
    shiftRegs_addressIn_delay_234_1 <= shiftRegs_addressIn_delay_233_1;
    shiftRegs_addressIn_delay_235_0 <= shiftRegs_addressIn_delay_234_0;
    shiftRegs_addressIn_delay_235_1 <= shiftRegs_addressIn_delay_234_1;
    shiftRegs_addressIn_delay_236_0 <= shiftRegs_addressIn_delay_235_0;
    shiftRegs_addressIn_delay_236_1 <= shiftRegs_addressIn_delay_235_1;
    shiftRegs_addressIn_delay_237_0 <= shiftRegs_addressIn_delay_236_0;
    shiftRegs_addressIn_delay_237_1 <= shiftRegs_addressIn_delay_236_1;
    shiftRegs_addressIn_delay_238_0 <= shiftRegs_addressIn_delay_237_0;
    shiftRegs_addressIn_delay_238_1 <= shiftRegs_addressIn_delay_237_1;
    shiftRegs_addressIn_delay_239_0 <= shiftRegs_addressIn_delay_238_0;
    shiftRegs_addressIn_delay_239_1 <= shiftRegs_addressIn_delay_238_1;
    shiftRegs_addressIn_delay_240_0 <= shiftRegs_addressIn_delay_239_0;
    shiftRegs_addressIn_delay_240_1 <= shiftRegs_addressIn_delay_239_1;
    shiftRegs_addressIn_delay_241_0 <= shiftRegs_addressIn_delay_240_0;
    shiftRegs_addressIn_delay_241_1 <= shiftRegs_addressIn_delay_240_1;
    shiftRegs_addressIn_delay_242_0 <= shiftRegs_addressIn_delay_241_0;
    shiftRegs_addressIn_delay_242_1 <= shiftRegs_addressIn_delay_241_1;
    shiftRegs_addressIn_delay_243_0 <= shiftRegs_addressIn_delay_242_0;
    shiftRegs_addressIn_delay_243_1 <= shiftRegs_addressIn_delay_242_1;
    shiftRegs_addressIn_delay_244_0 <= shiftRegs_addressIn_delay_243_0;
    shiftRegs_addressIn_delay_244_1 <= shiftRegs_addressIn_delay_243_1;
    shiftRegs_addressIn_delay_245_0 <= shiftRegs_addressIn_delay_244_0;
    shiftRegs_addressIn_delay_245_1 <= shiftRegs_addressIn_delay_244_1;
    shiftRegs_addressIn_delay_246_0 <= shiftRegs_addressIn_delay_245_0;
    shiftRegs_addressIn_delay_246_1 <= shiftRegs_addressIn_delay_245_1;
    shiftRegs_addressIn_delay_247_0 <= shiftRegs_addressIn_delay_246_0;
    shiftRegs_addressIn_delay_247_1 <= shiftRegs_addressIn_delay_246_1;
    shiftRegs_addressIn_delay_248_0 <= shiftRegs_addressIn_delay_247_0;
    shiftRegs_addressIn_delay_248_1 <= shiftRegs_addressIn_delay_247_1;
    shiftRegs_addressIn_delay_249_0 <= shiftRegs_addressIn_delay_248_0;
    shiftRegs_addressIn_delay_249_1 <= shiftRegs_addressIn_delay_248_1;
    shiftRegs_addressIn_delay_250_0 <= shiftRegs_addressIn_delay_249_0;
    shiftRegs_addressIn_delay_250_1 <= shiftRegs_addressIn_delay_249_1;
    shiftRegs_addressIn_delay_251_0 <= shiftRegs_addressIn_delay_250_0;
    shiftRegs_addressIn_delay_251_1 <= shiftRegs_addressIn_delay_250_1;
    shiftRegs_addressIn_delay_252_0 <= shiftRegs_addressIn_delay_251_0;
    shiftRegs_addressIn_delay_252_1 <= shiftRegs_addressIn_delay_251_1;
    shiftRegs_addressIn_delay_253_0 <= shiftRegs_addressIn_delay_252_0;
    shiftRegs_addressIn_delay_253_1 <= shiftRegs_addressIn_delay_252_1;
    shiftRegs_addressIn_delay_254_0 <= shiftRegs_addressIn_delay_253_0;
    shiftRegs_addressIn_delay_254_1 <= shiftRegs_addressIn_delay_253_1;
    shiftRegs_addressOut_0 <= shiftRegs_addressIn_delay_254_0;
    shiftRegs_addressOut_1 <= shiftRegs_addressIn_delay_254_1;
    shiftRegs_addressOut_delay_1_0 <= shiftRegs_addressOut_0;
    shiftRegs_addressOut_delay_1_1 <= shiftRegs_addressOut_1;
    shiftRegs_addressOut_delay_2_0 <= shiftRegs_addressOut_delay_1_0;
    shiftRegs_addressOut_delay_2_1 <= shiftRegs_addressOut_delay_1_1;
    shiftRegs_addressOut_delay_3_0 <= shiftRegs_addressOut_delay_2_0;
    shiftRegs_addressOut_delay_3_1 <= shiftRegs_addressOut_delay_2_1;
    shiftRegs_addressOut_delay_4_0 <= shiftRegs_addressOut_delay_3_0;
    shiftRegs_addressOut_delay_4_1 <= shiftRegs_addressOut_delay_3_1;
    shiftRegs_addressOutFull_0 <= shiftRegs_addressOut_delay_4_0;
    shiftRegs_addressOutFull_1 <= shiftRegs_addressOut_delay_4_1;
    pAddPort_0_s_regNext_X <= pAddPort_0_s_X;
    pAddPort_0_s_regNext_Y <= pAddPort_0_s_Y;
    pAddPort_0_s_regNext_Z <= pAddPort_0_s_Z;
    pAddPort_0_s_regNext_T <= pAddPort_0_s_T;
    _zz_stage1_inputAddress_0 <= {stage1_GCnt_value,stage1_inputBarrelIDAbs_0};
    _zz_stage1_inputAddress_0_1 <= _zz_stage1_inputAddress_0;
    _zz_stage1_inputAddress_0_2 <= _zz_stage1_inputAddress_0_1;
    _zz_stage1_inputAddress_0_3 <= _zz_stage1_inputAddress_0_2;
    _zz_stage1_inputAddress_0_4 <= _zz_stage1_inputAddress_0_3;
    stage1_inputAddress_0 <= _zz_stage1_inputAddress_0_4;
    _zz_stage1_inputAddress_1 <= {stage1_GCnt_value,stage1_inputBarrelIDAbs_1};
    _zz_stage1_inputAddress_1_1 <= _zz_stage1_inputAddress_1;
    _zz_stage1_inputAddress_1_2 <= _zz_stage1_inputAddress_1_1;
    _zz_stage1_inputAddress_1_3 <= _zz_stage1_inputAddress_1_2;
    _zz_stage1_inputAddress_1_4 <= _zz_stage1_inputAddress_1_3;
    stage1_inputAddress_1 <= _zz_stage1_inputAddress_1_4;
    _zz_stage1_inputData_0_X <= stage1_inputBarrelID_0[12];
    _zz_stage1_inputData_0_X_1 <= _zz_stage1_inputData_0_X;
    _zz_stage1_inputData_0_X_2 <= _zz_stage1_inputData_0_X_1;
    _zz_stage1_inputData_0_X_3 <= _zz_stage1_inputData_0_X_2;
    _zz_stage1_inputData_0_X_4 <= _zz_stage1_inputData_0_X_3;
    _zz_stage1_inputData_0_X_5 <= _zz_stage1_inputData_0_X_4;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_X <= dataInBuffer_bufferOut_payload_fragment_P_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y <= dataInBuffer_bufferOut_payload_fragment_P_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z <= dataInBuffer_bufferOut_payload_fragment_P_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_T <= dataInBuffer_bufferOut_payload_fragment_P_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_T;
    _zz_stage1_inputData_1_X <= stage1_inputBarrelID_1[12];
    _zz_stage1_inputData_1_X_1 <= _zz_stage1_inputData_1_X;
    _zz_stage1_inputData_1_X_2 <= _zz_stage1_inputData_1_X_1;
    _zz_stage1_inputData_1_X_3 <= _zz_stage1_inputData_1_X_2;
    _zz_stage1_inputData_1_X_4 <= _zz_stage1_inputData_1_X_3;
    _zz_stage1_inputData_1_X_5 <= _zz_stage1_inputData_1_X_4;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_X_1 <= dataInBuffer_bufferOut_payload_fragment_P_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y_1 <= dataInBuffer_bufferOut_payload_fragment_P_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z_1 <= dataInBuffer_bufferOut_payload_fragment_P_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_T_1 <= dataInBuffer_bufferOut_payload_fragment_P_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_X_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_X_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_T_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_T_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_X_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_X_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_T_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_T_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_X_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_X_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_T_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_T_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_X_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_X_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_T_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_T_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_X_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_X_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z_1;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_T_1 <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_T_1;
  end

  always @(posedge clk) begin
    stage1_inputValid_0_delay_1 <= stage1_inputValid_0;
    stage1_inputValid_0_delay_2 <= stage1_inputValid_0_delay_1;
    stage1_inputValid_0_delay_3 <= stage1_inputValid_0_delay_2;
    stage1_inputValid_0_delay_4 <= stage1_inputValid_0_delay_3;
    stage1_inputValid_0_delay_5 <= stage1_inputValid_0_delay_4;
    stage1_inputAddress_0_delay_1 <= stage1_inputAddress_0;
    stage1_inputAddress_0_delay_2 <= stage1_inputAddress_0_delay_1;
    stage1_inputAddress_0_delay_3 <= stage1_inputAddress_0_delay_2;
    stage1_inputAddress_0_delay_4 <= stage1_inputAddress_0_delay_3;
    stage1_inputAddress_0_delay_5 <= stage1_inputAddress_0_delay_4;
    stage1_inputData_0_delay_1_X <= stage1_inputData_0_X;
    stage1_inputData_0_delay_1_Y <= stage1_inputData_0_Y;
    stage1_inputData_0_delay_1_Z <= stage1_inputData_0_Z;
    stage1_inputData_0_delay_1_T <= stage1_inputData_0_T;
    stage1_inputData_0_delay_2_X <= stage1_inputData_0_delay_1_X;
    stage1_inputData_0_delay_2_Y <= stage1_inputData_0_delay_1_Y;
    stage1_inputData_0_delay_2_Z <= stage1_inputData_0_delay_1_Z;
    stage1_inputData_0_delay_2_T <= stage1_inputData_0_delay_1_T;
    stage1_inputData_0_delay_3_X <= stage1_inputData_0_delay_2_X;
    stage1_inputData_0_delay_3_Y <= stage1_inputData_0_delay_2_Y;
    stage1_inputData_0_delay_3_Z <= stage1_inputData_0_delay_2_Z;
    stage1_inputData_0_delay_3_T <= stage1_inputData_0_delay_2_T;
    stage1_inputData_0_delay_4_X <= stage1_inputData_0_delay_3_X;
    stage1_inputData_0_delay_4_Y <= stage1_inputData_0_delay_3_Y;
    stage1_inputData_0_delay_4_Z <= stage1_inputData_0_delay_3_Z;
    stage1_inputData_0_delay_4_T <= stage1_inputData_0_delay_3_T;
    stage1_inputData_0_delay_5_X <= stage1_inputData_0_delay_4_X;
    stage1_inputData_0_delay_5_Y <= stage1_inputData_0_delay_4_Y;
    stage1_inputData_0_delay_5_Z <= stage1_inputData_0_delay_4_Z;
    stage1_inputData_0_delay_5_T <= stage1_inputData_0_delay_4_T;
    _zz_io_dataIn_0_valid <= (stage1_inputValid_0 && (stage1_inputAddress_0 == shiftRegs_addressOut_0));
    _zz_io_dataIn_0_valid_1 <= _zz_io_dataIn_0_valid;
    _zz_io_dataIn_0_valid_2 <= _zz_io_dataIn_0_valid_1;
    _zz_io_dataIn_0_valid_3 <= _zz_io_dataIn_0_valid_2;
    _zz_io_dataIn_0_valid_4 <= _zz_io_dataIn_0_valid_3;
    _zz_io_dataIn_0_payload_a_X <= (stage1_inputValid_0 && (stage1_inputAddress_0 == shiftRegs_addressOut_0));
    _zz_io_dataIn_0_payload_a_X_1 <= _zz_io_dataIn_0_payload_a_X;
    _zz_io_dataIn_0_payload_a_X_2 <= _zz_io_dataIn_0_payload_a_X_1;
    _zz_io_dataIn_0_payload_a_X_3 <= _zz_io_dataIn_0_payload_a_X_2;
    _zz_io_dataIn_0_payload_a_X_4 <= _zz_io_dataIn_0_payload_a_X_3;
    _zz_io_dataIn_0_payload_a_X_5 <= _zz_io_dataIn_0_payload_a_X_4;
    _zz_io_dataIn_0_payload_a_X_6 <= _zz_io_dataIn_0_payload_a_X_5;
    _zz_io_dataIn_0_payload_a_X_7 <= _zz_io_dataIn_0_payload_a_X_6;
    _zz_io_dataIn_0_payload_a_X_8 <= _zz_io_dataIn_0_payload_a_X_7;
    _zz_io_dataIn_0_payload_a_X_9 <= _zz_io_dataIn_0_payload_a_X_8;
    _zz_io_dataIn_0_payload_a_X_10 <= _zz_io_dataIn_0_payload_a_X_9;
    _zz_io_dataIn_0_payload_a_X_11 <= _zz_io_dataIn_0_payload_a_X_10;
    _zz_io_dataIn_0_payload_a_X_12 <= _zz_io_dataIn_0_payload_a_X_11;
    _zz_io_dataIn_0_payload_a_X_13 <= _zz_io_dataIn_0_payload_a_X_12;
    _zz_io_dataIn_0_payload_a_X_14 <= _zz_io_dataIn_0_payload_a_X_13;
    _zz_io_dataIn_0_payload_a_X_15 <= _zz_io_dataIn_0_payload_a_X_14;
    _zz_io_dataIn_0_payload_a_X_16 <= _zz_io_dataIn_0_payload_a_X_15;
    _zz_io_dataIn_0_payload_a_X_17 <= _zz_io_dataIn_0_payload_a_X_16;
    _zz_io_dataIn_0_payload_a_X_18 <= _zz_io_dataIn_0_payload_a_X_17;
    _zz_io_dataIn_0_payload_a_X_19 <= _zz_io_dataIn_0_payload_a_X_18;
    _zz_io_dataIn_0_payload_a_X_20 <= _zz_io_dataIn_0_payload_a_X_19;
    _zz_io_dataIn_0_payload_a_X_21 <= _zz_io_dataIn_0_payload_a_X_20;
    _zz_io_dataIn_0_payload_a_X_22 <= _zz_io_dataIn_0_payload_a_X_21;
    _zz_io_dataIn_0_payload_a_X_23 <= _zz_io_dataIn_0_payload_a_X_22;
    _zz_io_dataIn_0_payload_a_X_24 <= _zz_io_dataIn_0_payload_a_X_23;
    _zz_io_dataIn_0_payload_a_X_25 <= _zz_io_dataIn_0_payload_a_X_24;
    _zz_io_dataIn_0_payload_a_X_26 <= _zz_io_dataIn_0_payload_a_X_25;
    _zz_io_dataIn_0_payload_a_X_27 <= _zz_io_dataIn_0_payload_a_X_26;
    _zz_io_dataIn_0_payload_a_X_28 <= _zz_io_dataIn_0_payload_a_X_27;
    _zz_io_dataIn_0_payload_a_X_29 <= _zz_io_dataIn_0_payload_a_X_28;
    _zz_io_dataIn_0_payload_a_X_30 <= _zz_io_dataIn_0_payload_a_X_29;
    _zz_io_dataIn_0_payload_a_X_31 <= _zz_io_dataIn_0_payload_a_X_30;
    _zz_io_dataIn_0_payload_a_X_32 <= _zz_io_dataIn_0_payload_a_X_31;
    _zz_io_dataIn_0_payload_a_X_33 <= _zz_io_dataIn_0_payload_a_X_32;
    _zz_io_dataIn_0_payload_a_X_34 <= _zz_io_dataIn_0_payload_a_X_33;
    stage1_inputData_0_delay_1_X_1 <= stage1_inputData_0_X;
    stage1_inputData_0_delay_1_Y_1 <= stage1_inputData_0_Y;
    stage1_inputData_0_delay_1_Z_1 <= stage1_inputData_0_Z;
    stage1_inputData_0_delay_1_T_1 <= stage1_inputData_0_T;
    stage1_inputData_0_delay_2_X_1 <= stage1_inputData_0_delay_1_X_1;
    stage1_inputData_0_delay_2_Y_1 <= stage1_inputData_0_delay_1_Y_1;
    stage1_inputData_0_delay_2_Z_1 <= stage1_inputData_0_delay_1_Z_1;
    stage1_inputData_0_delay_2_T_1 <= stage1_inputData_0_delay_1_T_1;
    stage1_inputData_0_delay_3_X_1 <= stage1_inputData_0_delay_2_X_1;
    stage1_inputData_0_delay_3_Y_1 <= stage1_inputData_0_delay_2_Y_1;
    stage1_inputData_0_delay_3_Z_1 <= stage1_inputData_0_delay_2_Z_1;
    stage1_inputData_0_delay_3_T_1 <= stage1_inputData_0_delay_2_T_1;
    stage1_inputData_0_delay_4_X_1 <= stage1_inputData_0_delay_3_X_1;
    stage1_inputData_0_delay_4_Y_1 <= stage1_inputData_0_delay_3_Y_1;
    stage1_inputData_0_delay_4_Z_1 <= stage1_inputData_0_delay_3_Z_1;
    stage1_inputData_0_delay_4_T_1 <= stage1_inputData_0_delay_3_T_1;
    stage1_inputData_0_delay_5_X_1 <= stage1_inputData_0_delay_4_X_1;
    stage1_inputData_0_delay_5_Y_1 <= stage1_inputData_0_delay_4_Y_1;
    stage1_inputData_0_delay_5_Z_1 <= stage1_inputData_0_delay_4_Z_1;
    stage1_inputData_0_delay_5_T_1 <= stage1_inputData_0_delay_4_T_1;
    stage1_inputData_0_delay_6_X <= stage1_inputData_0_delay_5_X_1;
    stage1_inputData_0_delay_6_Y <= stage1_inputData_0_delay_5_Y_1;
    stage1_inputData_0_delay_6_Z <= stage1_inputData_0_delay_5_Z_1;
    stage1_inputData_0_delay_6_T <= stage1_inputData_0_delay_5_T_1;
    stage1_inputData_0_delay_7_X <= stage1_inputData_0_delay_6_X;
    stage1_inputData_0_delay_7_Y <= stage1_inputData_0_delay_6_Y;
    stage1_inputData_0_delay_7_Z <= stage1_inputData_0_delay_6_Z;
    stage1_inputData_0_delay_7_T <= stage1_inputData_0_delay_6_T;
    stage1_inputData_0_delay_8_X <= stage1_inputData_0_delay_7_X;
    stage1_inputData_0_delay_8_Y <= stage1_inputData_0_delay_7_Y;
    stage1_inputData_0_delay_8_Z <= stage1_inputData_0_delay_7_Z;
    stage1_inputData_0_delay_8_T <= stage1_inputData_0_delay_7_T;
    stage1_inputData_0_delay_9_X <= stage1_inputData_0_delay_8_X;
    stage1_inputData_0_delay_9_Y <= stage1_inputData_0_delay_8_Y;
    stage1_inputData_0_delay_9_Z <= stage1_inputData_0_delay_8_Z;
    stage1_inputData_0_delay_9_T <= stage1_inputData_0_delay_8_T;
    stage1_inputData_0_delay_10_X <= stage1_inputData_0_delay_9_X;
    stage1_inputData_0_delay_10_Y <= stage1_inputData_0_delay_9_Y;
    stage1_inputData_0_delay_10_Z <= stage1_inputData_0_delay_9_Z;
    stage1_inputData_0_delay_10_T <= stage1_inputData_0_delay_9_T;
    stage1_inputData_0_delay_11_X <= stage1_inputData_0_delay_10_X;
    stage1_inputData_0_delay_11_Y <= stage1_inputData_0_delay_10_Y;
    stage1_inputData_0_delay_11_Z <= stage1_inputData_0_delay_10_Z;
    stage1_inputData_0_delay_11_T <= stage1_inputData_0_delay_10_T;
    stage1_inputData_0_delay_12_X <= stage1_inputData_0_delay_11_X;
    stage1_inputData_0_delay_12_Y <= stage1_inputData_0_delay_11_Y;
    stage1_inputData_0_delay_12_Z <= stage1_inputData_0_delay_11_Z;
    stage1_inputData_0_delay_12_T <= stage1_inputData_0_delay_11_T;
    stage1_inputData_0_delay_13_X <= stage1_inputData_0_delay_12_X;
    stage1_inputData_0_delay_13_Y <= stage1_inputData_0_delay_12_Y;
    stage1_inputData_0_delay_13_Z <= stage1_inputData_0_delay_12_Z;
    stage1_inputData_0_delay_13_T <= stage1_inputData_0_delay_12_T;
    stage1_inputData_0_delay_14_X <= stage1_inputData_0_delay_13_X;
    stage1_inputData_0_delay_14_Y <= stage1_inputData_0_delay_13_Y;
    stage1_inputData_0_delay_14_Z <= stage1_inputData_0_delay_13_Z;
    stage1_inputData_0_delay_14_T <= stage1_inputData_0_delay_13_T;
    stage1_inputData_0_delay_15_X <= stage1_inputData_0_delay_14_X;
    stage1_inputData_0_delay_15_Y <= stage1_inputData_0_delay_14_Y;
    stage1_inputData_0_delay_15_Z <= stage1_inputData_0_delay_14_Z;
    stage1_inputData_0_delay_15_T <= stage1_inputData_0_delay_14_T;
    stage1_inputData_0_delay_16_X <= stage1_inputData_0_delay_15_X;
    stage1_inputData_0_delay_16_Y <= stage1_inputData_0_delay_15_Y;
    stage1_inputData_0_delay_16_Z <= stage1_inputData_0_delay_15_Z;
    stage1_inputData_0_delay_16_T <= stage1_inputData_0_delay_15_T;
    stage1_inputData_0_delay_17_X <= stage1_inputData_0_delay_16_X;
    stage1_inputData_0_delay_17_Y <= stage1_inputData_0_delay_16_Y;
    stage1_inputData_0_delay_17_Z <= stage1_inputData_0_delay_16_Z;
    stage1_inputData_0_delay_17_T <= stage1_inputData_0_delay_16_T;
    stage1_inputData_0_delay_18_X <= stage1_inputData_0_delay_17_X;
    stage1_inputData_0_delay_18_Y <= stage1_inputData_0_delay_17_Y;
    stage1_inputData_0_delay_18_Z <= stage1_inputData_0_delay_17_Z;
    stage1_inputData_0_delay_18_T <= stage1_inputData_0_delay_17_T;
    stage1_inputData_0_delay_19_X <= stage1_inputData_0_delay_18_X;
    stage1_inputData_0_delay_19_Y <= stage1_inputData_0_delay_18_Y;
    stage1_inputData_0_delay_19_Z <= stage1_inputData_0_delay_18_Z;
    stage1_inputData_0_delay_19_T <= stage1_inputData_0_delay_18_T;
    stage1_inputData_0_delay_20_X <= stage1_inputData_0_delay_19_X;
    stage1_inputData_0_delay_20_Y <= stage1_inputData_0_delay_19_Y;
    stage1_inputData_0_delay_20_Z <= stage1_inputData_0_delay_19_Z;
    stage1_inputData_0_delay_20_T <= stage1_inputData_0_delay_19_T;
    stage1_inputData_0_delay_21_X <= stage1_inputData_0_delay_20_X;
    stage1_inputData_0_delay_21_Y <= stage1_inputData_0_delay_20_Y;
    stage1_inputData_0_delay_21_Z <= stage1_inputData_0_delay_20_Z;
    stage1_inputData_0_delay_21_T <= stage1_inputData_0_delay_20_T;
    stage1_inputData_0_delay_22_X <= stage1_inputData_0_delay_21_X;
    stage1_inputData_0_delay_22_Y <= stage1_inputData_0_delay_21_Y;
    stage1_inputData_0_delay_22_Z <= stage1_inputData_0_delay_21_Z;
    stage1_inputData_0_delay_22_T <= stage1_inputData_0_delay_21_T;
    stage1_inputData_0_delay_23_X <= stage1_inputData_0_delay_22_X;
    stage1_inputData_0_delay_23_Y <= stage1_inputData_0_delay_22_Y;
    stage1_inputData_0_delay_23_Z <= stage1_inputData_0_delay_22_Z;
    stage1_inputData_0_delay_23_T <= stage1_inputData_0_delay_22_T;
    stage1_inputData_0_delay_24_X <= stage1_inputData_0_delay_23_X;
    stage1_inputData_0_delay_24_Y <= stage1_inputData_0_delay_23_Y;
    stage1_inputData_0_delay_24_Z <= stage1_inputData_0_delay_23_Z;
    stage1_inputData_0_delay_24_T <= stage1_inputData_0_delay_23_T;
    stage1_inputData_0_delay_25_X <= stage1_inputData_0_delay_24_X;
    stage1_inputData_0_delay_25_Y <= stage1_inputData_0_delay_24_Y;
    stage1_inputData_0_delay_25_Z <= stage1_inputData_0_delay_24_Z;
    stage1_inputData_0_delay_25_T <= stage1_inputData_0_delay_24_T;
    stage1_inputData_0_delay_26_X <= stage1_inputData_0_delay_25_X;
    stage1_inputData_0_delay_26_Y <= stage1_inputData_0_delay_25_Y;
    stage1_inputData_0_delay_26_Z <= stage1_inputData_0_delay_25_Z;
    stage1_inputData_0_delay_26_T <= stage1_inputData_0_delay_25_T;
    stage1_inputData_0_delay_27_X <= stage1_inputData_0_delay_26_X;
    stage1_inputData_0_delay_27_Y <= stage1_inputData_0_delay_26_Y;
    stage1_inputData_0_delay_27_Z <= stage1_inputData_0_delay_26_Z;
    stage1_inputData_0_delay_27_T <= stage1_inputData_0_delay_26_T;
    stage1_inputData_0_delay_28_X <= stage1_inputData_0_delay_27_X;
    stage1_inputData_0_delay_28_Y <= stage1_inputData_0_delay_27_Y;
    stage1_inputData_0_delay_28_Z <= stage1_inputData_0_delay_27_Z;
    stage1_inputData_0_delay_28_T <= stage1_inputData_0_delay_27_T;
    stage1_inputData_0_delay_29_X <= stage1_inputData_0_delay_28_X;
    stage1_inputData_0_delay_29_Y <= stage1_inputData_0_delay_28_Y;
    stage1_inputData_0_delay_29_Z <= stage1_inputData_0_delay_28_Z;
    stage1_inputData_0_delay_29_T <= stage1_inputData_0_delay_28_T;
    stage1_inputData_0_delay_30_X <= stage1_inputData_0_delay_29_X;
    stage1_inputData_0_delay_30_Y <= stage1_inputData_0_delay_29_Y;
    stage1_inputData_0_delay_30_Z <= stage1_inputData_0_delay_29_Z;
    stage1_inputData_0_delay_30_T <= stage1_inputData_0_delay_29_T;
    stage1_inputData_0_delay_31_X <= stage1_inputData_0_delay_30_X;
    stage1_inputData_0_delay_31_Y <= stage1_inputData_0_delay_30_Y;
    stage1_inputData_0_delay_31_Z <= stage1_inputData_0_delay_30_Z;
    stage1_inputData_0_delay_31_T <= stage1_inputData_0_delay_30_T;
    stage1_inputData_0_delay_32_X <= stage1_inputData_0_delay_31_X;
    stage1_inputData_0_delay_32_Y <= stage1_inputData_0_delay_31_Y;
    stage1_inputData_0_delay_32_Z <= stage1_inputData_0_delay_31_Z;
    stage1_inputData_0_delay_32_T <= stage1_inputData_0_delay_31_T;
    stage1_inputData_0_delay_33_X <= stage1_inputData_0_delay_32_X;
    stage1_inputData_0_delay_33_Y <= stage1_inputData_0_delay_32_Y;
    stage1_inputData_0_delay_33_Z <= stage1_inputData_0_delay_32_Z;
    stage1_inputData_0_delay_33_T <= stage1_inputData_0_delay_32_T;
    stage1_inputData_0_delay_34_X <= stage1_inputData_0_delay_33_X;
    stage1_inputData_0_delay_34_Y <= stage1_inputData_0_delay_33_Y;
    stage1_inputData_0_delay_34_Z <= stage1_inputData_0_delay_33_Z;
    stage1_inputData_0_delay_34_T <= stage1_inputData_0_delay_33_T;
    stage1_inputData_0_delay_35_X <= stage1_inputData_0_delay_34_X;
    stage1_inputData_0_delay_35_Y <= stage1_inputData_0_delay_34_Y;
    stage1_inputData_0_delay_35_Z <= stage1_inputData_0_delay_34_Z;
    stage1_inputData_0_delay_35_T <= stage1_inputData_0_delay_34_T;
    pAddPort_0_s_delay_1_X <= pAddPort_0_s_X;
    pAddPort_0_s_delay_1_Y <= pAddPort_0_s_Y;
    pAddPort_0_s_delay_1_Z <= pAddPort_0_s_Z;
    pAddPort_0_s_delay_1_T <= pAddPort_0_s_T;
    pAddPort_0_s_delay_2_X <= pAddPort_0_s_delay_1_X;
    pAddPort_0_s_delay_2_Y <= pAddPort_0_s_delay_1_Y;
    pAddPort_0_s_delay_2_Z <= pAddPort_0_s_delay_1_Z;
    pAddPort_0_s_delay_2_T <= pAddPort_0_s_delay_1_T;
    pAddPort_0_s_delay_3_X <= pAddPort_0_s_delay_2_X;
    pAddPort_0_s_delay_3_Y <= pAddPort_0_s_delay_2_Y;
    pAddPort_0_s_delay_3_Z <= pAddPort_0_s_delay_2_Z;
    pAddPort_0_s_delay_3_T <= pAddPort_0_s_delay_2_T;
    pAddPort_0_s_delay_4_X <= pAddPort_0_s_delay_3_X;
    pAddPort_0_s_delay_4_Y <= pAddPort_0_s_delay_3_Y;
    pAddPort_0_s_delay_4_Z <= pAddPort_0_s_delay_3_Z;
    pAddPort_0_s_delay_4_T <= pAddPort_0_s_delay_3_T;
    pAddPort_0_s_delay_5_X <= pAddPort_0_s_delay_4_X;
    pAddPort_0_s_delay_5_Y <= pAddPort_0_s_delay_4_Y;
    pAddPort_0_s_delay_5_Z <= pAddPort_0_s_delay_4_Z;
    pAddPort_0_s_delay_5_T <= pAddPort_0_s_delay_4_T;
    pAddPort_0_s_delay_6_X <= pAddPort_0_s_delay_5_X;
    pAddPort_0_s_delay_6_Y <= pAddPort_0_s_delay_5_Y;
    pAddPort_0_s_delay_6_Z <= pAddPort_0_s_delay_5_Z;
    pAddPort_0_s_delay_6_T <= pAddPort_0_s_delay_5_T;
    pAddPort_0_s_delay_7_X <= pAddPort_0_s_delay_6_X;
    pAddPort_0_s_delay_7_Y <= pAddPort_0_s_delay_6_Y;
    pAddPort_0_s_delay_7_Z <= pAddPort_0_s_delay_6_Z;
    pAddPort_0_s_delay_7_T <= pAddPort_0_s_delay_6_T;
    pAddPort_0_s_delay_8_X <= pAddPort_0_s_delay_7_X;
    pAddPort_0_s_delay_8_Y <= pAddPort_0_s_delay_7_Y;
    pAddPort_0_s_delay_8_Z <= pAddPort_0_s_delay_7_Z;
    pAddPort_0_s_delay_8_T <= pAddPort_0_s_delay_7_T;
    pAddPort_0_s_delay_9_X <= pAddPort_0_s_delay_8_X;
    pAddPort_0_s_delay_9_Y <= pAddPort_0_s_delay_8_Y;
    pAddPort_0_s_delay_9_Z <= pAddPort_0_s_delay_8_Z;
    pAddPort_0_s_delay_9_T <= pAddPort_0_s_delay_8_T;
    pAddPort_0_s_delay_10_X <= pAddPort_0_s_delay_9_X;
    pAddPort_0_s_delay_10_Y <= pAddPort_0_s_delay_9_Y;
    pAddPort_0_s_delay_10_Z <= pAddPort_0_s_delay_9_Z;
    pAddPort_0_s_delay_10_T <= pAddPort_0_s_delay_9_T;
    pAddPort_0_s_delay_11_X <= pAddPort_0_s_delay_10_X;
    pAddPort_0_s_delay_11_Y <= pAddPort_0_s_delay_10_Y;
    pAddPort_0_s_delay_11_Z <= pAddPort_0_s_delay_10_Z;
    pAddPort_0_s_delay_11_T <= pAddPort_0_s_delay_10_T;
    pAddPort_0_s_delay_12_X <= pAddPort_0_s_delay_11_X;
    pAddPort_0_s_delay_12_Y <= pAddPort_0_s_delay_11_Y;
    pAddPort_0_s_delay_12_Z <= pAddPort_0_s_delay_11_Z;
    pAddPort_0_s_delay_12_T <= pAddPort_0_s_delay_11_T;
    pAddPort_0_s_delay_13_X <= pAddPort_0_s_delay_12_X;
    pAddPort_0_s_delay_13_Y <= pAddPort_0_s_delay_12_Y;
    pAddPort_0_s_delay_13_Z <= pAddPort_0_s_delay_12_Z;
    pAddPort_0_s_delay_13_T <= pAddPort_0_s_delay_12_T;
    pAddPort_0_s_delay_14_X <= pAddPort_0_s_delay_13_X;
    pAddPort_0_s_delay_14_Y <= pAddPort_0_s_delay_13_Y;
    pAddPort_0_s_delay_14_Z <= pAddPort_0_s_delay_13_Z;
    pAddPort_0_s_delay_14_T <= pAddPort_0_s_delay_13_T;
    pAddPort_0_s_delay_15_X <= pAddPort_0_s_delay_14_X;
    pAddPort_0_s_delay_15_Y <= pAddPort_0_s_delay_14_Y;
    pAddPort_0_s_delay_15_Z <= pAddPort_0_s_delay_14_Z;
    pAddPort_0_s_delay_15_T <= pAddPort_0_s_delay_14_T;
    pAddPort_0_s_delay_16_X <= pAddPort_0_s_delay_15_X;
    pAddPort_0_s_delay_16_Y <= pAddPort_0_s_delay_15_Y;
    pAddPort_0_s_delay_16_Z <= pAddPort_0_s_delay_15_Z;
    pAddPort_0_s_delay_16_T <= pAddPort_0_s_delay_15_T;
    pAddPort_0_s_delay_17_X <= pAddPort_0_s_delay_16_X;
    pAddPort_0_s_delay_17_Y <= pAddPort_0_s_delay_16_Y;
    pAddPort_0_s_delay_17_Z <= pAddPort_0_s_delay_16_Z;
    pAddPort_0_s_delay_17_T <= pAddPort_0_s_delay_16_T;
    pAddPort_0_s_delay_18_X <= pAddPort_0_s_delay_17_X;
    pAddPort_0_s_delay_18_Y <= pAddPort_0_s_delay_17_Y;
    pAddPort_0_s_delay_18_Z <= pAddPort_0_s_delay_17_Z;
    pAddPort_0_s_delay_18_T <= pAddPort_0_s_delay_17_T;
    pAddPort_0_s_delay_19_X <= pAddPort_0_s_delay_18_X;
    pAddPort_0_s_delay_19_Y <= pAddPort_0_s_delay_18_Y;
    pAddPort_0_s_delay_19_Z <= pAddPort_0_s_delay_18_Z;
    pAddPort_0_s_delay_19_T <= pAddPort_0_s_delay_18_T;
    pAddPort_0_s_delay_20_X <= pAddPort_0_s_delay_19_X;
    pAddPort_0_s_delay_20_Y <= pAddPort_0_s_delay_19_Y;
    pAddPort_0_s_delay_20_Z <= pAddPort_0_s_delay_19_Z;
    pAddPort_0_s_delay_20_T <= pAddPort_0_s_delay_19_T;
    pAddPort_0_s_delay_21_X <= pAddPort_0_s_delay_20_X;
    pAddPort_0_s_delay_21_Y <= pAddPort_0_s_delay_20_Y;
    pAddPort_0_s_delay_21_Z <= pAddPort_0_s_delay_20_Z;
    pAddPort_0_s_delay_21_T <= pAddPort_0_s_delay_20_T;
    pAddPort_0_s_delay_22_X <= pAddPort_0_s_delay_21_X;
    pAddPort_0_s_delay_22_Y <= pAddPort_0_s_delay_21_Y;
    pAddPort_0_s_delay_22_Z <= pAddPort_0_s_delay_21_Z;
    pAddPort_0_s_delay_22_T <= pAddPort_0_s_delay_21_T;
    pAddPort_0_s_delay_23_X <= pAddPort_0_s_delay_22_X;
    pAddPort_0_s_delay_23_Y <= pAddPort_0_s_delay_22_Y;
    pAddPort_0_s_delay_23_Z <= pAddPort_0_s_delay_22_Z;
    pAddPort_0_s_delay_23_T <= pAddPort_0_s_delay_22_T;
    pAddPort_0_s_delay_24_X <= pAddPort_0_s_delay_23_X;
    pAddPort_0_s_delay_24_Y <= pAddPort_0_s_delay_23_Y;
    pAddPort_0_s_delay_24_Z <= pAddPort_0_s_delay_23_Z;
    pAddPort_0_s_delay_24_T <= pAddPort_0_s_delay_23_T;
    pAddPort_0_s_delay_25_X <= pAddPort_0_s_delay_24_X;
    pAddPort_0_s_delay_25_Y <= pAddPort_0_s_delay_24_Y;
    pAddPort_0_s_delay_25_Z <= pAddPort_0_s_delay_24_Z;
    pAddPort_0_s_delay_25_T <= pAddPort_0_s_delay_24_T;
    pAddPort_0_s_delay_26_X <= pAddPort_0_s_delay_25_X;
    pAddPort_0_s_delay_26_Y <= pAddPort_0_s_delay_25_Y;
    pAddPort_0_s_delay_26_Z <= pAddPort_0_s_delay_25_Z;
    pAddPort_0_s_delay_26_T <= pAddPort_0_s_delay_25_T;
    pAddPort_0_s_delay_27_X <= pAddPort_0_s_delay_26_X;
    pAddPort_0_s_delay_27_Y <= pAddPort_0_s_delay_26_Y;
    pAddPort_0_s_delay_27_Z <= pAddPort_0_s_delay_26_Z;
    pAddPort_0_s_delay_27_T <= pAddPort_0_s_delay_26_T;
    pAddPort_0_s_delay_28_X <= pAddPort_0_s_delay_27_X;
    pAddPort_0_s_delay_28_Y <= pAddPort_0_s_delay_27_Y;
    pAddPort_0_s_delay_28_Z <= pAddPort_0_s_delay_27_Z;
    pAddPort_0_s_delay_28_T <= pAddPort_0_s_delay_27_T;
    pAddPort_0_s_delay_29_X <= pAddPort_0_s_delay_28_X;
    pAddPort_0_s_delay_29_Y <= pAddPort_0_s_delay_28_Y;
    pAddPort_0_s_delay_29_Z <= pAddPort_0_s_delay_28_Z;
    pAddPort_0_s_delay_29_T <= pAddPort_0_s_delay_28_T;
    pAddPort_0_s_delay_30_X <= pAddPort_0_s_delay_29_X;
    pAddPort_0_s_delay_30_Y <= pAddPort_0_s_delay_29_Y;
    pAddPort_0_s_delay_30_Z <= pAddPort_0_s_delay_29_Z;
    pAddPort_0_s_delay_30_T <= pAddPort_0_s_delay_29_T;
    shiftRegs_addressOutFull_0_delay_1 <= shiftRegs_addressOutFull_0;
    shiftRegs_addressOutFull_0_delay_2 <= shiftRegs_addressOutFull_0_delay_1;
    shiftRegs_addressOutFull_0_delay_3 <= shiftRegs_addressOutFull_0_delay_2;
    shiftRegs_addressOutFull_0_delay_4 <= shiftRegs_addressOutFull_0_delay_3;
    shiftRegs_addressOutFull_0_delay_5 <= shiftRegs_addressOutFull_0_delay_4;
    shiftRegs_addressOutFull_0_delay_6 <= shiftRegs_addressOutFull_0_delay_5;
    shiftRegs_addressOutFull_0_delay_7 <= shiftRegs_addressOutFull_0_delay_6;
    shiftRegs_addressOutFull_0_delay_8 <= shiftRegs_addressOutFull_0_delay_7;
    shiftRegs_addressOutFull_0_delay_9 <= shiftRegs_addressOutFull_0_delay_8;
    shiftRegs_addressOutFull_0_delay_10 <= shiftRegs_addressOutFull_0_delay_9;
    shiftRegs_addressOutFull_0_delay_11 <= shiftRegs_addressOutFull_0_delay_10;
    shiftRegs_addressOutFull_0_delay_12 <= shiftRegs_addressOutFull_0_delay_11;
    shiftRegs_addressOutFull_0_delay_13 <= shiftRegs_addressOutFull_0_delay_12;
    shiftRegs_addressOutFull_0_delay_14 <= shiftRegs_addressOutFull_0_delay_13;
    shiftRegs_addressOutFull_0_delay_15 <= shiftRegs_addressOutFull_0_delay_14;
    shiftRegs_addressOutFull_0_delay_16 <= shiftRegs_addressOutFull_0_delay_15;
    shiftRegs_addressOutFull_0_delay_17 <= shiftRegs_addressOutFull_0_delay_16;
    shiftRegs_addressOutFull_0_delay_18 <= shiftRegs_addressOutFull_0_delay_17;
    shiftRegs_addressOutFull_0_delay_19 <= shiftRegs_addressOutFull_0_delay_18;
    shiftRegs_addressOutFull_0_delay_20 <= shiftRegs_addressOutFull_0_delay_19;
    shiftRegs_addressOutFull_0_delay_21 <= shiftRegs_addressOutFull_0_delay_20;
    shiftRegs_addressOutFull_0_delay_22 <= shiftRegs_addressOutFull_0_delay_21;
    shiftRegs_addressOutFull_0_delay_23 <= shiftRegs_addressOutFull_0_delay_22;
    shiftRegs_addressOutFull_0_delay_24 <= shiftRegs_addressOutFull_0_delay_23;
    shiftRegs_addressOutFull_0_delay_25 <= shiftRegs_addressOutFull_0_delay_24;
    shiftRegs_addressOutFull_0_delay_26 <= shiftRegs_addressOutFull_0_delay_25;
    shiftRegs_addressOutFull_0_delay_27 <= shiftRegs_addressOutFull_0_delay_26;
    shiftRegs_addressOutFull_0_delay_28 <= shiftRegs_addressOutFull_0_delay_27;
    shiftRegs_addressOutFull_0_delay_29 <= shiftRegs_addressOutFull_0_delay_28;
    shiftRegs_addressOutFull_0_delay_30 <= shiftRegs_addressOutFull_0_delay_29;
    stage1_inputData_0_delay_1_X_2 <= stage1_inputData_0_X;
    stage1_inputData_0_delay_1_Y_2 <= stage1_inputData_0_Y;
    stage1_inputData_0_delay_1_Z_2 <= stage1_inputData_0_Z;
    stage1_inputData_0_delay_1_T_2 <= stage1_inputData_0_T;
    stage1_inputData_0_delay_2_X_2 <= stage1_inputData_0_delay_1_X_2;
    stage1_inputData_0_delay_2_Y_2 <= stage1_inputData_0_delay_1_Y_2;
    stage1_inputData_0_delay_2_Z_2 <= stage1_inputData_0_delay_1_Z_2;
    stage1_inputData_0_delay_2_T_2 <= stage1_inputData_0_delay_1_T_2;
    stage1_inputData_0_delay_3_X_2 <= stage1_inputData_0_delay_2_X_2;
    stage1_inputData_0_delay_3_Y_2 <= stage1_inputData_0_delay_2_Y_2;
    stage1_inputData_0_delay_3_Z_2 <= stage1_inputData_0_delay_2_Z_2;
    stage1_inputData_0_delay_3_T_2 <= stage1_inputData_0_delay_2_T_2;
    stage1_inputData_0_delay_4_X_2 <= stage1_inputData_0_delay_3_X_2;
    stage1_inputData_0_delay_4_Y_2 <= stage1_inputData_0_delay_3_Y_2;
    stage1_inputData_0_delay_4_Z_2 <= stage1_inputData_0_delay_3_Z_2;
    stage1_inputData_0_delay_4_T_2 <= stage1_inputData_0_delay_3_T_2;
    stage1_inputData_0_delay_5_X_2 <= stage1_inputData_0_delay_4_X_2;
    stage1_inputData_0_delay_5_Y_2 <= stage1_inputData_0_delay_4_Y_2;
    stage1_inputData_0_delay_5_Z_2 <= stage1_inputData_0_delay_4_Z_2;
    stage1_inputData_0_delay_5_T_2 <= stage1_inputData_0_delay_4_T_2;
    stage1_inputData_0_delay_6_X_1 <= stage1_inputData_0_delay_5_X_2;
    stage1_inputData_0_delay_6_Y_1 <= stage1_inputData_0_delay_5_Y_2;
    stage1_inputData_0_delay_6_Z_1 <= stage1_inputData_0_delay_5_Z_2;
    stage1_inputData_0_delay_6_T_1 <= stage1_inputData_0_delay_5_T_2;
    stage1_inputData_0_delay_7_X_1 <= stage1_inputData_0_delay_6_X_1;
    stage1_inputData_0_delay_7_Y_1 <= stage1_inputData_0_delay_6_Y_1;
    stage1_inputData_0_delay_7_Z_1 <= stage1_inputData_0_delay_6_Z_1;
    stage1_inputData_0_delay_7_T_1 <= stage1_inputData_0_delay_6_T_1;
    stage1_inputData_0_delay_8_X_1 <= stage1_inputData_0_delay_7_X_1;
    stage1_inputData_0_delay_8_Y_1 <= stage1_inputData_0_delay_7_Y_1;
    stage1_inputData_0_delay_8_Z_1 <= stage1_inputData_0_delay_7_Z_1;
    stage1_inputData_0_delay_8_T_1 <= stage1_inputData_0_delay_7_T_1;
    stage1_inputData_0_delay_9_X_1 <= stage1_inputData_0_delay_8_X_1;
    stage1_inputData_0_delay_9_Y_1 <= stage1_inputData_0_delay_8_Y_1;
    stage1_inputData_0_delay_9_Z_1 <= stage1_inputData_0_delay_8_Z_1;
    stage1_inputData_0_delay_9_T_1 <= stage1_inputData_0_delay_8_T_1;
    stage1_inputData_0_delay_10_X_1 <= stage1_inputData_0_delay_9_X_1;
    stage1_inputData_0_delay_10_Y_1 <= stage1_inputData_0_delay_9_Y_1;
    stage1_inputData_0_delay_10_Z_1 <= stage1_inputData_0_delay_9_Z_1;
    stage1_inputData_0_delay_10_T_1 <= stage1_inputData_0_delay_9_T_1;
    stage1_inputData_0_delay_11_X_1 <= stage1_inputData_0_delay_10_X_1;
    stage1_inputData_0_delay_11_Y_1 <= stage1_inputData_0_delay_10_Y_1;
    stage1_inputData_0_delay_11_Z_1 <= stage1_inputData_0_delay_10_Z_1;
    stage1_inputData_0_delay_11_T_1 <= stage1_inputData_0_delay_10_T_1;
    stage1_inputData_0_delay_12_X_1 <= stage1_inputData_0_delay_11_X_1;
    stage1_inputData_0_delay_12_Y_1 <= stage1_inputData_0_delay_11_Y_1;
    stage1_inputData_0_delay_12_Z_1 <= stage1_inputData_0_delay_11_Z_1;
    stage1_inputData_0_delay_12_T_1 <= stage1_inputData_0_delay_11_T_1;
    stage1_inputData_0_delay_13_X_1 <= stage1_inputData_0_delay_12_X_1;
    stage1_inputData_0_delay_13_Y_1 <= stage1_inputData_0_delay_12_Y_1;
    stage1_inputData_0_delay_13_Z_1 <= stage1_inputData_0_delay_12_Z_1;
    stage1_inputData_0_delay_13_T_1 <= stage1_inputData_0_delay_12_T_1;
    stage1_inputData_0_delay_14_X_1 <= stage1_inputData_0_delay_13_X_1;
    stage1_inputData_0_delay_14_Y_1 <= stage1_inputData_0_delay_13_Y_1;
    stage1_inputData_0_delay_14_Z_1 <= stage1_inputData_0_delay_13_Z_1;
    stage1_inputData_0_delay_14_T_1 <= stage1_inputData_0_delay_13_T_1;
    stage1_inputData_0_delay_15_X_1 <= stage1_inputData_0_delay_14_X_1;
    stage1_inputData_0_delay_15_Y_1 <= stage1_inputData_0_delay_14_Y_1;
    stage1_inputData_0_delay_15_Z_1 <= stage1_inputData_0_delay_14_Z_1;
    stage1_inputData_0_delay_15_T_1 <= stage1_inputData_0_delay_14_T_1;
    stage1_inputData_0_delay_16_X_1 <= stage1_inputData_0_delay_15_X_1;
    stage1_inputData_0_delay_16_Y_1 <= stage1_inputData_0_delay_15_Y_1;
    stage1_inputData_0_delay_16_Z_1 <= stage1_inputData_0_delay_15_Z_1;
    stage1_inputData_0_delay_16_T_1 <= stage1_inputData_0_delay_15_T_1;
    stage1_inputData_0_delay_17_X_1 <= stage1_inputData_0_delay_16_X_1;
    stage1_inputData_0_delay_17_Y_1 <= stage1_inputData_0_delay_16_Y_1;
    stage1_inputData_0_delay_17_Z_1 <= stage1_inputData_0_delay_16_Z_1;
    stage1_inputData_0_delay_17_T_1 <= stage1_inputData_0_delay_16_T_1;
    stage1_inputData_0_delay_18_X_1 <= stage1_inputData_0_delay_17_X_1;
    stage1_inputData_0_delay_18_Y_1 <= stage1_inputData_0_delay_17_Y_1;
    stage1_inputData_0_delay_18_Z_1 <= stage1_inputData_0_delay_17_Z_1;
    stage1_inputData_0_delay_18_T_1 <= stage1_inputData_0_delay_17_T_1;
    stage1_inputData_0_delay_19_X_1 <= stage1_inputData_0_delay_18_X_1;
    stage1_inputData_0_delay_19_Y_1 <= stage1_inputData_0_delay_18_Y_1;
    stage1_inputData_0_delay_19_Z_1 <= stage1_inputData_0_delay_18_Z_1;
    stage1_inputData_0_delay_19_T_1 <= stage1_inputData_0_delay_18_T_1;
    stage1_inputData_0_delay_20_X_1 <= stage1_inputData_0_delay_19_X_1;
    stage1_inputData_0_delay_20_Y_1 <= stage1_inputData_0_delay_19_Y_1;
    stage1_inputData_0_delay_20_Z_1 <= stage1_inputData_0_delay_19_Z_1;
    stage1_inputData_0_delay_20_T_1 <= stage1_inputData_0_delay_19_T_1;
    stage1_inputData_0_delay_21_X_1 <= stage1_inputData_0_delay_20_X_1;
    stage1_inputData_0_delay_21_Y_1 <= stage1_inputData_0_delay_20_Y_1;
    stage1_inputData_0_delay_21_Z_1 <= stage1_inputData_0_delay_20_Z_1;
    stage1_inputData_0_delay_21_T_1 <= stage1_inputData_0_delay_20_T_1;
    stage1_inputData_0_delay_22_X_1 <= stage1_inputData_0_delay_21_X_1;
    stage1_inputData_0_delay_22_Y_1 <= stage1_inputData_0_delay_21_Y_1;
    stage1_inputData_0_delay_22_Z_1 <= stage1_inputData_0_delay_21_Z_1;
    stage1_inputData_0_delay_22_T_1 <= stage1_inputData_0_delay_21_T_1;
    stage1_inputData_0_delay_23_X_1 <= stage1_inputData_0_delay_22_X_1;
    stage1_inputData_0_delay_23_Y_1 <= stage1_inputData_0_delay_22_Y_1;
    stage1_inputData_0_delay_23_Z_1 <= stage1_inputData_0_delay_22_Z_1;
    stage1_inputData_0_delay_23_T_1 <= stage1_inputData_0_delay_22_T_1;
    stage1_inputData_0_delay_24_X_1 <= stage1_inputData_0_delay_23_X_1;
    stage1_inputData_0_delay_24_Y_1 <= stage1_inputData_0_delay_23_Y_1;
    stage1_inputData_0_delay_24_Z_1 <= stage1_inputData_0_delay_23_Z_1;
    stage1_inputData_0_delay_24_T_1 <= stage1_inputData_0_delay_23_T_1;
    stage1_inputData_0_delay_25_X_1 <= stage1_inputData_0_delay_24_X_1;
    stage1_inputData_0_delay_25_Y_1 <= stage1_inputData_0_delay_24_Y_1;
    stage1_inputData_0_delay_25_Z_1 <= stage1_inputData_0_delay_24_Z_1;
    stage1_inputData_0_delay_25_T_1 <= stage1_inputData_0_delay_24_T_1;
    stage1_inputData_0_delay_26_X_1 <= stage1_inputData_0_delay_25_X_1;
    stage1_inputData_0_delay_26_Y_1 <= stage1_inputData_0_delay_25_Y_1;
    stage1_inputData_0_delay_26_Z_1 <= stage1_inputData_0_delay_25_Z_1;
    stage1_inputData_0_delay_26_T_1 <= stage1_inputData_0_delay_25_T_1;
    stage1_inputData_0_delay_27_X_1 <= stage1_inputData_0_delay_26_X_1;
    stage1_inputData_0_delay_27_Y_1 <= stage1_inputData_0_delay_26_Y_1;
    stage1_inputData_0_delay_27_Z_1 <= stage1_inputData_0_delay_26_Z_1;
    stage1_inputData_0_delay_27_T_1 <= stage1_inputData_0_delay_26_T_1;
    stage1_inputData_0_delay_28_X_1 <= stage1_inputData_0_delay_27_X_1;
    stage1_inputData_0_delay_28_Y_1 <= stage1_inputData_0_delay_27_Y_1;
    stage1_inputData_0_delay_28_Z_1 <= stage1_inputData_0_delay_27_Z_1;
    stage1_inputData_0_delay_28_T_1 <= stage1_inputData_0_delay_27_T_1;
    stage1_inputData_0_delay_29_X_1 <= stage1_inputData_0_delay_28_X_1;
    stage1_inputData_0_delay_29_Y_1 <= stage1_inputData_0_delay_28_Y_1;
    stage1_inputData_0_delay_29_Z_1 <= stage1_inputData_0_delay_28_Z_1;
    stage1_inputData_0_delay_29_T_1 <= stage1_inputData_0_delay_28_T_1;
    stage1_inputData_0_delay_30_X_1 <= stage1_inputData_0_delay_29_X_1;
    stage1_inputData_0_delay_30_Y_1 <= stage1_inputData_0_delay_29_Y_1;
    stage1_inputData_0_delay_30_Z_1 <= stage1_inputData_0_delay_29_Z_1;
    stage1_inputData_0_delay_30_T_1 <= stage1_inputData_0_delay_29_T_1;
    stage1_inputData_0_delay_31_X_1 <= stage1_inputData_0_delay_30_X_1;
    stage1_inputData_0_delay_31_Y_1 <= stage1_inputData_0_delay_30_Y_1;
    stage1_inputData_0_delay_31_Z_1 <= stage1_inputData_0_delay_30_Z_1;
    stage1_inputData_0_delay_31_T_1 <= stage1_inputData_0_delay_30_T_1;
    stage1_inputData_0_delay_32_X_1 <= stage1_inputData_0_delay_31_X_1;
    stage1_inputData_0_delay_32_Y_1 <= stage1_inputData_0_delay_31_Y_1;
    stage1_inputData_0_delay_32_Z_1 <= stage1_inputData_0_delay_31_Z_1;
    stage1_inputData_0_delay_32_T_1 <= stage1_inputData_0_delay_31_T_1;
    stage1_inputData_0_delay_33_X_1 <= stage1_inputData_0_delay_32_X_1;
    stage1_inputData_0_delay_33_Y_1 <= stage1_inputData_0_delay_32_Y_1;
    stage1_inputData_0_delay_33_Z_1 <= stage1_inputData_0_delay_32_Z_1;
    stage1_inputData_0_delay_33_T_1 <= stage1_inputData_0_delay_32_T_1;
    stage1_inputData_0_delay_34_X_1 <= stage1_inputData_0_delay_33_X_1;
    stage1_inputData_0_delay_34_Y_1 <= stage1_inputData_0_delay_33_Y_1;
    stage1_inputData_0_delay_34_Z_1 <= stage1_inputData_0_delay_33_Z_1;
    stage1_inputData_0_delay_34_T_1 <= stage1_inputData_0_delay_33_T_1;
    stage1_inputData_0_delay_35_X_1 <= stage1_inputData_0_delay_34_X_1;
    stage1_inputData_0_delay_35_Y_1 <= stage1_inputData_0_delay_34_Y_1;
    stage1_inputData_0_delay_35_Z_1 <= stage1_inputData_0_delay_34_Z_1;
    stage1_inputData_0_delay_35_T_1 <= stage1_inputData_0_delay_34_T_1;
    stage1_inputAddress_0_delay_1_1 <= stage1_inputAddress_0;
    stage1_inputAddress_0_delay_2_1 <= stage1_inputAddress_0_delay_1_1;
    stage1_inputAddress_0_delay_3_1 <= stage1_inputAddress_0_delay_2_1;
    stage1_inputAddress_0_delay_4_1 <= stage1_inputAddress_0_delay_3_1;
    stage1_inputAddress_0_delay_5_1 <= stage1_inputAddress_0_delay_4_1;
    stage1_inputAddress_0_delay_6 <= stage1_inputAddress_0_delay_5_1;
    stage1_inputAddress_0_delay_7 <= stage1_inputAddress_0_delay_6;
    stage1_inputAddress_0_delay_8 <= stage1_inputAddress_0_delay_7;
    stage1_inputAddress_0_delay_9 <= stage1_inputAddress_0_delay_8;
    stage1_inputAddress_0_delay_10 <= stage1_inputAddress_0_delay_9;
    stage1_inputAddress_0_delay_11 <= stage1_inputAddress_0_delay_10;
    stage1_inputAddress_0_delay_12 <= stage1_inputAddress_0_delay_11;
    stage1_inputAddress_0_delay_13 <= stage1_inputAddress_0_delay_12;
    stage1_inputAddress_0_delay_14 <= stage1_inputAddress_0_delay_13;
    stage1_inputAddress_0_delay_15 <= stage1_inputAddress_0_delay_14;
    stage1_inputAddress_0_delay_16 <= stage1_inputAddress_0_delay_15;
    stage1_inputAddress_0_delay_17 <= stage1_inputAddress_0_delay_16;
    stage1_inputAddress_0_delay_18 <= stage1_inputAddress_0_delay_17;
    stage1_inputAddress_0_delay_19 <= stage1_inputAddress_0_delay_18;
    stage1_inputAddress_0_delay_20 <= stage1_inputAddress_0_delay_19;
    stage1_inputAddress_0_delay_21 <= stage1_inputAddress_0_delay_20;
    stage1_inputAddress_0_delay_22 <= stage1_inputAddress_0_delay_21;
    stage1_inputAddress_0_delay_23 <= stage1_inputAddress_0_delay_22;
    stage1_inputAddress_0_delay_24 <= stage1_inputAddress_0_delay_23;
    stage1_inputAddress_0_delay_25 <= stage1_inputAddress_0_delay_24;
    stage1_inputAddress_0_delay_26 <= stage1_inputAddress_0_delay_25;
    stage1_inputAddress_0_delay_27 <= stage1_inputAddress_0_delay_26;
    stage1_inputAddress_0_delay_28 <= stage1_inputAddress_0_delay_27;
    stage1_inputAddress_0_delay_29 <= stage1_inputAddress_0_delay_28;
    stage1_inputAddress_0_delay_30 <= stage1_inputAddress_0_delay_29;
    stage1_inputAddress_0_delay_31 <= stage1_inputAddress_0_delay_30;
    stage1_inputAddress_0_delay_32 <= stage1_inputAddress_0_delay_31;
    stage1_inputAddress_0_delay_33 <= stage1_inputAddress_0_delay_32;
    stage1_inputAddress_0_delay_34 <= stage1_inputAddress_0_delay_33;
    stage1_inputAddress_0_delay_35 <= stage1_inputAddress_0_delay_34;
    stage1_inputValid_1_delay_1 <= stage1_inputValid_1;
    stage1_inputValid_1_delay_2 <= stage1_inputValid_1_delay_1;
    stage1_inputValid_1_delay_3 <= stage1_inputValid_1_delay_2;
    stage1_inputValid_1_delay_4 <= stage1_inputValid_1_delay_3;
    stage1_inputValid_1_delay_5 <= stage1_inputValid_1_delay_4;
    stage1_inputAddress_1_delay_1 <= stage1_inputAddress_1;
    stage1_inputAddress_1_delay_2 <= stage1_inputAddress_1_delay_1;
    stage1_inputAddress_1_delay_3 <= stage1_inputAddress_1_delay_2;
    stage1_inputAddress_1_delay_4 <= stage1_inputAddress_1_delay_3;
    stage1_inputAddress_1_delay_5 <= stage1_inputAddress_1_delay_4;
    stage1_inputData_1_delay_1_X <= stage1_inputData_1_X;
    stage1_inputData_1_delay_1_Y <= stage1_inputData_1_Y;
    stage1_inputData_1_delay_1_Z <= stage1_inputData_1_Z;
    stage1_inputData_1_delay_1_T <= stage1_inputData_1_T;
    stage1_inputData_1_delay_2_X <= stage1_inputData_1_delay_1_X;
    stage1_inputData_1_delay_2_Y <= stage1_inputData_1_delay_1_Y;
    stage1_inputData_1_delay_2_Z <= stage1_inputData_1_delay_1_Z;
    stage1_inputData_1_delay_2_T <= stage1_inputData_1_delay_1_T;
    stage1_inputData_1_delay_3_X <= stage1_inputData_1_delay_2_X;
    stage1_inputData_1_delay_3_Y <= stage1_inputData_1_delay_2_Y;
    stage1_inputData_1_delay_3_Z <= stage1_inputData_1_delay_2_Z;
    stage1_inputData_1_delay_3_T <= stage1_inputData_1_delay_2_T;
    stage1_inputData_1_delay_4_X <= stage1_inputData_1_delay_3_X;
    stage1_inputData_1_delay_4_Y <= stage1_inputData_1_delay_3_Y;
    stage1_inputData_1_delay_4_Z <= stage1_inputData_1_delay_3_Z;
    stage1_inputData_1_delay_4_T <= stage1_inputData_1_delay_3_T;
    stage1_inputData_1_delay_5_X <= stage1_inputData_1_delay_4_X;
    stage1_inputData_1_delay_5_Y <= stage1_inputData_1_delay_4_Y;
    stage1_inputData_1_delay_5_Z <= stage1_inputData_1_delay_4_Z;
    stage1_inputData_1_delay_5_T <= stage1_inputData_1_delay_4_T;
    _zz_io_dataIn_0_valid_35 <= (stage1_inputValid_1 && (stage1_inputAddress_1 == shiftRegs_addressOut_1));
    _zz_io_dataIn_0_valid_36 <= _zz_io_dataIn_0_valid_35;
    _zz_io_dataIn_0_valid_37 <= _zz_io_dataIn_0_valid_36;
    _zz_io_dataIn_0_valid_38 <= _zz_io_dataIn_0_valid_37;
    _zz_io_dataIn_0_valid_39 <= _zz_io_dataIn_0_valid_38;
    _zz_io_dataIn_0_payload_a_X_35 <= (stage1_inputValid_1 && (stage1_inputAddress_1 == shiftRegs_addressOut_1));
    _zz_io_dataIn_0_payload_a_X_36 <= _zz_io_dataIn_0_payload_a_X_35;
    _zz_io_dataIn_0_payload_a_X_37 <= _zz_io_dataIn_0_payload_a_X_36;
    _zz_io_dataIn_0_payload_a_X_38 <= _zz_io_dataIn_0_payload_a_X_37;
    _zz_io_dataIn_0_payload_a_X_39 <= _zz_io_dataIn_0_payload_a_X_38;
    _zz_io_dataIn_0_payload_a_X_40 <= _zz_io_dataIn_0_payload_a_X_39;
    _zz_io_dataIn_0_payload_a_X_41 <= _zz_io_dataIn_0_payload_a_X_40;
    _zz_io_dataIn_0_payload_a_X_42 <= _zz_io_dataIn_0_payload_a_X_41;
    _zz_io_dataIn_0_payload_a_X_43 <= _zz_io_dataIn_0_payload_a_X_42;
    _zz_io_dataIn_0_payload_a_X_44 <= _zz_io_dataIn_0_payload_a_X_43;
    _zz_io_dataIn_0_payload_a_X_45 <= _zz_io_dataIn_0_payload_a_X_44;
    _zz_io_dataIn_0_payload_a_X_46 <= _zz_io_dataIn_0_payload_a_X_45;
    _zz_io_dataIn_0_payload_a_X_47 <= _zz_io_dataIn_0_payload_a_X_46;
    _zz_io_dataIn_0_payload_a_X_48 <= _zz_io_dataIn_0_payload_a_X_47;
    _zz_io_dataIn_0_payload_a_X_49 <= _zz_io_dataIn_0_payload_a_X_48;
    _zz_io_dataIn_0_payload_a_X_50 <= _zz_io_dataIn_0_payload_a_X_49;
    _zz_io_dataIn_0_payload_a_X_51 <= _zz_io_dataIn_0_payload_a_X_50;
    _zz_io_dataIn_0_payload_a_X_52 <= _zz_io_dataIn_0_payload_a_X_51;
    _zz_io_dataIn_0_payload_a_X_53 <= _zz_io_dataIn_0_payload_a_X_52;
    _zz_io_dataIn_0_payload_a_X_54 <= _zz_io_dataIn_0_payload_a_X_53;
    _zz_io_dataIn_0_payload_a_X_55 <= _zz_io_dataIn_0_payload_a_X_54;
    _zz_io_dataIn_0_payload_a_X_56 <= _zz_io_dataIn_0_payload_a_X_55;
    _zz_io_dataIn_0_payload_a_X_57 <= _zz_io_dataIn_0_payload_a_X_56;
    _zz_io_dataIn_0_payload_a_X_58 <= _zz_io_dataIn_0_payload_a_X_57;
    _zz_io_dataIn_0_payload_a_X_59 <= _zz_io_dataIn_0_payload_a_X_58;
    _zz_io_dataIn_0_payload_a_X_60 <= _zz_io_dataIn_0_payload_a_X_59;
    _zz_io_dataIn_0_payload_a_X_61 <= _zz_io_dataIn_0_payload_a_X_60;
    _zz_io_dataIn_0_payload_a_X_62 <= _zz_io_dataIn_0_payload_a_X_61;
    _zz_io_dataIn_0_payload_a_X_63 <= _zz_io_dataIn_0_payload_a_X_62;
    _zz_io_dataIn_0_payload_a_X_64 <= _zz_io_dataIn_0_payload_a_X_63;
    _zz_io_dataIn_0_payload_a_X_65 <= _zz_io_dataIn_0_payload_a_X_64;
    _zz_io_dataIn_0_payload_a_X_66 <= _zz_io_dataIn_0_payload_a_X_65;
    _zz_io_dataIn_0_payload_a_X_67 <= _zz_io_dataIn_0_payload_a_X_66;
    _zz_io_dataIn_0_payload_a_X_68 <= _zz_io_dataIn_0_payload_a_X_67;
    _zz_io_dataIn_0_payload_a_X_69 <= _zz_io_dataIn_0_payload_a_X_68;
    stage1_inputData_1_delay_1_X_1 <= stage1_inputData_1_X;
    stage1_inputData_1_delay_1_Y_1 <= stage1_inputData_1_Y;
    stage1_inputData_1_delay_1_Z_1 <= stage1_inputData_1_Z;
    stage1_inputData_1_delay_1_T_1 <= stage1_inputData_1_T;
    stage1_inputData_1_delay_2_X_1 <= stage1_inputData_1_delay_1_X_1;
    stage1_inputData_1_delay_2_Y_1 <= stage1_inputData_1_delay_1_Y_1;
    stage1_inputData_1_delay_2_Z_1 <= stage1_inputData_1_delay_1_Z_1;
    stage1_inputData_1_delay_2_T_1 <= stage1_inputData_1_delay_1_T_1;
    stage1_inputData_1_delay_3_X_1 <= stage1_inputData_1_delay_2_X_1;
    stage1_inputData_1_delay_3_Y_1 <= stage1_inputData_1_delay_2_Y_1;
    stage1_inputData_1_delay_3_Z_1 <= stage1_inputData_1_delay_2_Z_1;
    stage1_inputData_1_delay_3_T_1 <= stage1_inputData_1_delay_2_T_1;
    stage1_inputData_1_delay_4_X_1 <= stage1_inputData_1_delay_3_X_1;
    stage1_inputData_1_delay_4_Y_1 <= stage1_inputData_1_delay_3_Y_1;
    stage1_inputData_1_delay_4_Z_1 <= stage1_inputData_1_delay_3_Z_1;
    stage1_inputData_1_delay_4_T_1 <= stage1_inputData_1_delay_3_T_1;
    stage1_inputData_1_delay_5_X_1 <= stage1_inputData_1_delay_4_X_1;
    stage1_inputData_1_delay_5_Y_1 <= stage1_inputData_1_delay_4_Y_1;
    stage1_inputData_1_delay_5_Z_1 <= stage1_inputData_1_delay_4_Z_1;
    stage1_inputData_1_delay_5_T_1 <= stage1_inputData_1_delay_4_T_1;
    stage1_inputData_1_delay_6_X <= stage1_inputData_1_delay_5_X_1;
    stage1_inputData_1_delay_6_Y <= stage1_inputData_1_delay_5_Y_1;
    stage1_inputData_1_delay_6_Z <= stage1_inputData_1_delay_5_Z_1;
    stage1_inputData_1_delay_6_T <= stage1_inputData_1_delay_5_T_1;
    stage1_inputData_1_delay_7_X <= stage1_inputData_1_delay_6_X;
    stage1_inputData_1_delay_7_Y <= stage1_inputData_1_delay_6_Y;
    stage1_inputData_1_delay_7_Z <= stage1_inputData_1_delay_6_Z;
    stage1_inputData_1_delay_7_T <= stage1_inputData_1_delay_6_T;
    stage1_inputData_1_delay_8_X <= stage1_inputData_1_delay_7_X;
    stage1_inputData_1_delay_8_Y <= stage1_inputData_1_delay_7_Y;
    stage1_inputData_1_delay_8_Z <= stage1_inputData_1_delay_7_Z;
    stage1_inputData_1_delay_8_T <= stage1_inputData_1_delay_7_T;
    stage1_inputData_1_delay_9_X <= stage1_inputData_1_delay_8_X;
    stage1_inputData_1_delay_9_Y <= stage1_inputData_1_delay_8_Y;
    stage1_inputData_1_delay_9_Z <= stage1_inputData_1_delay_8_Z;
    stage1_inputData_1_delay_9_T <= stage1_inputData_1_delay_8_T;
    stage1_inputData_1_delay_10_X <= stage1_inputData_1_delay_9_X;
    stage1_inputData_1_delay_10_Y <= stage1_inputData_1_delay_9_Y;
    stage1_inputData_1_delay_10_Z <= stage1_inputData_1_delay_9_Z;
    stage1_inputData_1_delay_10_T <= stage1_inputData_1_delay_9_T;
    stage1_inputData_1_delay_11_X <= stage1_inputData_1_delay_10_X;
    stage1_inputData_1_delay_11_Y <= stage1_inputData_1_delay_10_Y;
    stage1_inputData_1_delay_11_Z <= stage1_inputData_1_delay_10_Z;
    stage1_inputData_1_delay_11_T <= stage1_inputData_1_delay_10_T;
    stage1_inputData_1_delay_12_X <= stage1_inputData_1_delay_11_X;
    stage1_inputData_1_delay_12_Y <= stage1_inputData_1_delay_11_Y;
    stage1_inputData_1_delay_12_Z <= stage1_inputData_1_delay_11_Z;
    stage1_inputData_1_delay_12_T <= stage1_inputData_1_delay_11_T;
    stage1_inputData_1_delay_13_X <= stage1_inputData_1_delay_12_X;
    stage1_inputData_1_delay_13_Y <= stage1_inputData_1_delay_12_Y;
    stage1_inputData_1_delay_13_Z <= stage1_inputData_1_delay_12_Z;
    stage1_inputData_1_delay_13_T <= stage1_inputData_1_delay_12_T;
    stage1_inputData_1_delay_14_X <= stage1_inputData_1_delay_13_X;
    stage1_inputData_1_delay_14_Y <= stage1_inputData_1_delay_13_Y;
    stage1_inputData_1_delay_14_Z <= stage1_inputData_1_delay_13_Z;
    stage1_inputData_1_delay_14_T <= stage1_inputData_1_delay_13_T;
    stage1_inputData_1_delay_15_X <= stage1_inputData_1_delay_14_X;
    stage1_inputData_1_delay_15_Y <= stage1_inputData_1_delay_14_Y;
    stage1_inputData_1_delay_15_Z <= stage1_inputData_1_delay_14_Z;
    stage1_inputData_1_delay_15_T <= stage1_inputData_1_delay_14_T;
    stage1_inputData_1_delay_16_X <= stage1_inputData_1_delay_15_X;
    stage1_inputData_1_delay_16_Y <= stage1_inputData_1_delay_15_Y;
    stage1_inputData_1_delay_16_Z <= stage1_inputData_1_delay_15_Z;
    stage1_inputData_1_delay_16_T <= stage1_inputData_1_delay_15_T;
    stage1_inputData_1_delay_17_X <= stage1_inputData_1_delay_16_X;
    stage1_inputData_1_delay_17_Y <= stage1_inputData_1_delay_16_Y;
    stage1_inputData_1_delay_17_Z <= stage1_inputData_1_delay_16_Z;
    stage1_inputData_1_delay_17_T <= stage1_inputData_1_delay_16_T;
    stage1_inputData_1_delay_18_X <= stage1_inputData_1_delay_17_X;
    stage1_inputData_1_delay_18_Y <= stage1_inputData_1_delay_17_Y;
    stage1_inputData_1_delay_18_Z <= stage1_inputData_1_delay_17_Z;
    stage1_inputData_1_delay_18_T <= stage1_inputData_1_delay_17_T;
    stage1_inputData_1_delay_19_X <= stage1_inputData_1_delay_18_X;
    stage1_inputData_1_delay_19_Y <= stage1_inputData_1_delay_18_Y;
    stage1_inputData_1_delay_19_Z <= stage1_inputData_1_delay_18_Z;
    stage1_inputData_1_delay_19_T <= stage1_inputData_1_delay_18_T;
    stage1_inputData_1_delay_20_X <= stage1_inputData_1_delay_19_X;
    stage1_inputData_1_delay_20_Y <= stage1_inputData_1_delay_19_Y;
    stage1_inputData_1_delay_20_Z <= stage1_inputData_1_delay_19_Z;
    stage1_inputData_1_delay_20_T <= stage1_inputData_1_delay_19_T;
    stage1_inputData_1_delay_21_X <= stage1_inputData_1_delay_20_X;
    stage1_inputData_1_delay_21_Y <= stage1_inputData_1_delay_20_Y;
    stage1_inputData_1_delay_21_Z <= stage1_inputData_1_delay_20_Z;
    stage1_inputData_1_delay_21_T <= stage1_inputData_1_delay_20_T;
    stage1_inputData_1_delay_22_X <= stage1_inputData_1_delay_21_X;
    stage1_inputData_1_delay_22_Y <= stage1_inputData_1_delay_21_Y;
    stage1_inputData_1_delay_22_Z <= stage1_inputData_1_delay_21_Z;
    stage1_inputData_1_delay_22_T <= stage1_inputData_1_delay_21_T;
    stage1_inputData_1_delay_23_X <= stage1_inputData_1_delay_22_X;
    stage1_inputData_1_delay_23_Y <= stage1_inputData_1_delay_22_Y;
    stage1_inputData_1_delay_23_Z <= stage1_inputData_1_delay_22_Z;
    stage1_inputData_1_delay_23_T <= stage1_inputData_1_delay_22_T;
    stage1_inputData_1_delay_24_X <= stage1_inputData_1_delay_23_X;
    stage1_inputData_1_delay_24_Y <= stage1_inputData_1_delay_23_Y;
    stage1_inputData_1_delay_24_Z <= stage1_inputData_1_delay_23_Z;
    stage1_inputData_1_delay_24_T <= stage1_inputData_1_delay_23_T;
    stage1_inputData_1_delay_25_X <= stage1_inputData_1_delay_24_X;
    stage1_inputData_1_delay_25_Y <= stage1_inputData_1_delay_24_Y;
    stage1_inputData_1_delay_25_Z <= stage1_inputData_1_delay_24_Z;
    stage1_inputData_1_delay_25_T <= stage1_inputData_1_delay_24_T;
    stage1_inputData_1_delay_26_X <= stage1_inputData_1_delay_25_X;
    stage1_inputData_1_delay_26_Y <= stage1_inputData_1_delay_25_Y;
    stage1_inputData_1_delay_26_Z <= stage1_inputData_1_delay_25_Z;
    stage1_inputData_1_delay_26_T <= stage1_inputData_1_delay_25_T;
    stage1_inputData_1_delay_27_X <= stage1_inputData_1_delay_26_X;
    stage1_inputData_1_delay_27_Y <= stage1_inputData_1_delay_26_Y;
    stage1_inputData_1_delay_27_Z <= stage1_inputData_1_delay_26_Z;
    stage1_inputData_1_delay_27_T <= stage1_inputData_1_delay_26_T;
    stage1_inputData_1_delay_28_X <= stage1_inputData_1_delay_27_X;
    stage1_inputData_1_delay_28_Y <= stage1_inputData_1_delay_27_Y;
    stage1_inputData_1_delay_28_Z <= stage1_inputData_1_delay_27_Z;
    stage1_inputData_1_delay_28_T <= stage1_inputData_1_delay_27_T;
    stage1_inputData_1_delay_29_X <= stage1_inputData_1_delay_28_X;
    stage1_inputData_1_delay_29_Y <= stage1_inputData_1_delay_28_Y;
    stage1_inputData_1_delay_29_Z <= stage1_inputData_1_delay_28_Z;
    stage1_inputData_1_delay_29_T <= stage1_inputData_1_delay_28_T;
    stage1_inputData_1_delay_30_X <= stage1_inputData_1_delay_29_X;
    stage1_inputData_1_delay_30_Y <= stage1_inputData_1_delay_29_Y;
    stage1_inputData_1_delay_30_Z <= stage1_inputData_1_delay_29_Z;
    stage1_inputData_1_delay_30_T <= stage1_inputData_1_delay_29_T;
    stage1_inputData_1_delay_31_X <= stage1_inputData_1_delay_30_X;
    stage1_inputData_1_delay_31_Y <= stage1_inputData_1_delay_30_Y;
    stage1_inputData_1_delay_31_Z <= stage1_inputData_1_delay_30_Z;
    stage1_inputData_1_delay_31_T <= stage1_inputData_1_delay_30_T;
    stage1_inputData_1_delay_32_X <= stage1_inputData_1_delay_31_X;
    stage1_inputData_1_delay_32_Y <= stage1_inputData_1_delay_31_Y;
    stage1_inputData_1_delay_32_Z <= stage1_inputData_1_delay_31_Z;
    stage1_inputData_1_delay_32_T <= stage1_inputData_1_delay_31_T;
    stage1_inputData_1_delay_33_X <= stage1_inputData_1_delay_32_X;
    stage1_inputData_1_delay_33_Y <= stage1_inputData_1_delay_32_Y;
    stage1_inputData_1_delay_33_Z <= stage1_inputData_1_delay_32_Z;
    stage1_inputData_1_delay_33_T <= stage1_inputData_1_delay_32_T;
    stage1_inputData_1_delay_34_X <= stage1_inputData_1_delay_33_X;
    stage1_inputData_1_delay_34_Y <= stage1_inputData_1_delay_33_Y;
    stage1_inputData_1_delay_34_Z <= stage1_inputData_1_delay_33_Z;
    stage1_inputData_1_delay_34_T <= stage1_inputData_1_delay_33_T;
    stage1_inputData_1_delay_35_X <= stage1_inputData_1_delay_34_X;
    stage1_inputData_1_delay_35_Y <= stage1_inputData_1_delay_34_Y;
    stage1_inputData_1_delay_35_Z <= stage1_inputData_1_delay_34_Z;
    stage1_inputData_1_delay_35_T <= stage1_inputData_1_delay_34_T;
    pAddPort_1_s_delay_1_X <= pAddPort_1_s_X;
    pAddPort_1_s_delay_1_Y <= pAddPort_1_s_Y;
    pAddPort_1_s_delay_1_Z <= pAddPort_1_s_Z;
    pAddPort_1_s_delay_1_T <= pAddPort_1_s_T;
    pAddPort_1_s_delay_2_X <= pAddPort_1_s_delay_1_X;
    pAddPort_1_s_delay_2_Y <= pAddPort_1_s_delay_1_Y;
    pAddPort_1_s_delay_2_Z <= pAddPort_1_s_delay_1_Z;
    pAddPort_1_s_delay_2_T <= pAddPort_1_s_delay_1_T;
    pAddPort_1_s_delay_3_X <= pAddPort_1_s_delay_2_X;
    pAddPort_1_s_delay_3_Y <= pAddPort_1_s_delay_2_Y;
    pAddPort_1_s_delay_3_Z <= pAddPort_1_s_delay_2_Z;
    pAddPort_1_s_delay_3_T <= pAddPort_1_s_delay_2_T;
    pAddPort_1_s_delay_4_X <= pAddPort_1_s_delay_3_X;
    pAddPort_1_s_delay_4_Y <= pAddPort_1_s_delay_3_Y;
    pAddPort_1_s_delay_4_Z <= pAddPort_1_s_delay_3_Z;
    pAddPort_1_s_delay_4_T <= pAddPort_1_s_delay_3_T;
    pAddPort_1_s_delay_5_X <= pAddPort_1_s_delay_4_X;
    pAddPort_1_s_delay_5_Y <= pAddPort_1_s_delay_4_Y;
    pAddPort_1_s_delay_5_Z <= pAddPort_1_s_delay_4_Z;
    pAddPort_1_s_delay_5_T <= pAddPort_1_s_delay_4_T;
    pAddPort_1_s_delay_6_X <= pAddPort_1_s_delay_5_X;
    pAddPort_1_s_delay_6_Y <= pAddPort_1_s_delay_5_Y;
    pAddPort_1_s_delay_6_Z <= pAddPort_1_s_delay_5_Z;
    pAddPort_1_s_delay_6_T <= pAddPort_1_s_delay_5_T;
    pAddPort_1_s_delay_7_X <= pAddPort_1_s_delay_6_X;
    pAddPort_1_s_delay_7_Y <= pAddPort_1_s_delay_6_Y;
    pAddPort_1_s_delay_7_Z <= pAddPort_1_s_delay_6_Z;
    pAddPort_1_s_delay_7_T <= pAddPort_1_s_delay_6_T;
    pAddPort_1_s_delay_8_X <= pAddPort_1_s_delay_7_X;
    pAddPort_1_s_delay_8_Y <= pAddPort_1_s_delay_7_Y;
    pAddPort_1_s_delay_8_Z <= pAddPort_1_s_delay_7_Z;
    pAddPort_1_s_delay_8_T <= pAddPort_1_s_delay_7_T;
    pAddPort_1_s_delay_9_X <= pAddPort_1_s_delay_8_X;
    pAddPort_1_s_delay_9_Y <= pAddPort_1_s_delay_8_Y;
    pAddPort_1_s_delay_9_Z <= pAddPort_1_s_delay_8_Z;
    pAddPort_1_s_delay_9_T <= pAddPort_1_s_delay_8_T;
    pAddPort_1_s_delay_10_X <= pAddPort_1_s_delay_9_X;
    pAddPort_1_s_delay_10_Y <= pAddPort_1_s_delay_9_Y;
    pAddPort_1_s_delay_10_Z <= pAddPort_1_s_delay_9_Z;
    pAddPort_1_s_delay_10_T <= pAddPort_1_s_delay_9_T;
    pAddPort_1_s_delay_11_X <= pAddPort_1_s_delay_10_X;
    pAddPort_1_s_delay_11_Y <= pAddPort_1_s_delay_10_Y;
    pAddPort_1_s_delay_11_Z <= pAddPort_1_s_delay_10_Z;
    pAddPort_1_s_delay_11_T <= pAddPort_1_s_delay_10_T;
    pAddPort_1_s_delay_12_X <= pAddPort_1_s_delay_11_X;
    pAddPort_1_s_delay_12_Y <= pAddPort_1_s_delay_11_Y;
    pAddPort_1_s_delay_12_Z <= pAddPort_1_s_delay_11_Z;
    pAddPort_1_s_delay_12_T <= pAddPort_1_s_delay_11_T;
    pAddPort_1_s_delay_13_X <= pAddPort_1_s_delay_12_X;
    pAddPort_1_s_delay_13_Y <= pAddPort_1_s_delay_12_Y;
    pAddPort_1_s_delay_13_Z <= pAddPort_1_s_delay_12_Z;
    pAddPort_1_s_delay_13_T <= pAddPort_1_s_delay_12_T;
    pAddPort_1_s_delay_14_X <= pAddPort_1_s_delay_13_X;
    pAddPort_1_s_delay_14_Y <= pAddPort_1_s_delay_13_Y;
    pAddPort_1_s_delay_14_Z <= pAddPort_1_s_delay_13_Z;
    pAddPort_1_s_delay_14_T <= pAddPort_1_s_delay_13_T;
    pAddPort_1_s_delay_15_X <= pAddPort_1_s_delay_14_X;
    pAddPort_1_s_delay_15_Y <= pAddPort_1_s_delay_14_Y;
    pAddPort_1_s_delay_15_Z <= pAddPort_1_s_delay_14_Z;
    pAddPort_1_s_delay_15_T <= pAddPort_1_s_delay_14_T;
    pAddPort_1_s_delay_16_X <= pAddPort_1_s_delay_15_X;
    pAddPort_1_s_delay_16_Y <= pAddPort_1_s_delay_15_Y;
    pAddPort_1_s_delay_16_Z <= pAddPort_1_s_delay_15_Z;
    pAddPort_1_s_delay_16_T <= pAddPort_1_s_delay_15_T;
    pAddPort_1_s_delay_17_X <= pAddPort_1_s_delay_16_X;
    pAddPort_1_s_delay_17_Y <= pAddPort_1_s_delay_16_Y;
    pAddPort_1_s_delay_17_Z <= pAddPort_1_s_delay_16_Z;
    pAddPort_1_s_delay_17_T <= pAddPort_1_s_delay_16_T;
    pAddPort_1_s_delay_18_X <= pAddPort_1_s_delay_17_X;
    pAddPort_1_s_delay_18_Y <= pAddPort_1_s_delay_17_Y;
    pAddPort_1_s_delay_18_Z <= pAddPort_1_s_delay_17_Z;
    pAddPort_1_s_delay_18_T <= pAddPort_1_s_delay_17_T;
    pAddPort_1_s_delay_19_X <= pAddPort_1_s_delay_18_X;
    pAddPort_1_s_delay_19_Y <= pAddPort_1_s_delay_18_Y;
    pAddPort_1_s_delay_19_Z <= pAddPort_1_s_delay_18_Z;
    pAddPort_1_s_delay_19_T <= pAddPort_1_s_delay_18_T;
    pAddPort_1_s_delay_20_X <= pAddPort_1_s_delay_19_X;
    pAddPort_1_s_delay_20_Y <= pAddPort_1_s_delay_19_Y;
    pAddPort_1_s_delay_20_Z <= pAddPort_1_s_delay_19_Z;
    pAddPort_1_s_delay_20_T <= pAddPort_1_s_delay_19_T;
    pAddPort_1_s_delay_21_X <= pAddPort_1_s_delay_20_X;
    pAddPort_1_s_delay_21_Y <= pAddPort_1_s_delay_20_Y;
    pAddPort_1_s_delay_21_Z <= pAddPort_1_s_delay_20_Z;
    pAddPort_1_s_delay_21_T <= pAddPort_1_s_delay_20_T;
    pAddPort_1_s_delay_22_X <= pAddPort_1_s_delay_21_X;
    pAddPort_1_s_delay_22_Y <= pAddPort_1_s_delay_21_Y;
    pAddPort_1_s_delay_22_Z <= pAddPort_1_s_delay_21_Z;
    pAddPort_1_s_delay_22_T <= pAddPort_1_s_delay_21_T;
    pAddPort_1_s_delay_23_X <= pAddPort_1_s_delay_22_X;
    pAddPort_1_s_delay_23_Y <= pAddPort_1_s_delay_22_Y;
    pAddPort_1_s_delay_23_Z <= pAddPort_1_s_delay_22_Z;
    pAddPort_1_s_delay_23_T <= pAddPort_1_s_delay_22_T;
    pAddPort_1_s_delay_24_X <= pAddPort_1_s_delay_23_X;
    pAddPort_1_s_delay_24_Y <= pAddPort_1_s_delay_23_Y;
    pAddPort_1_s_delay_24_Z <= pAddPort_1_s_delay_23_Z;
    pAddPort_1_s_delay_24_T <= pAddPort_1_s_delay_23_T;
    pAddPort_1_s_delay_25_X <= pAddPort_1_s_delay_24_X;
    pAddPort_1_s_delay_25_Y <= pAddPort_1_s_delay_24_Y;
    pAddPort_1_s_delay_25_Z <= pAddPort_1_s_delay_24_Z;
    pAddPort_1_s_delay_25_T <= pAddPort_1_s_delay_24_T;
    pAddPort_1_s_delay_26_X <= pAddPort_1_s_delay_25_X;
    pAddPort_1_s_delay_26_Y <= pAddPort_1_s_delay_25_Y;
    pAddPort_1_s_delay_26_Z <= pAddPort_1_s_delay_25_Z;
    pAddPort_1_s_delay_26_T <= pAddPort_1_s_delay_25_T;
    pAddPort_1_s_delay_27_X <= pAddPort_1_s_delay_26_X;
    pAddPort_1_s_delay_27_Y <= pAddPort_1_s_delay_26_Y;
    pAddPort_1_s_delay_27_Z <= pAddPort_1_s_delay_26_Z;
    pAddPort_1_s_delay_27_T <= pAddPort_1_s_delay_26_T;
    pAddPort_1_s_delay_28_X <= pAddPort_1_s_delay_27_X;
    pAddPort_1_s_delay_28_Y <= pAddPort_1_s_delay_27_Y;
    pAddPort_1_s_delay_28_Z <= pAddPort_1_s_delay_27_Z;
    pAddPort_1_s_delay_28_T <= pAddPort_1_s_delay_27_T;
    pAddPort_1_s_delay_29_X <= pAddPort_1_s_delay_28_X;
    pAddPort_1_s_delay_29_Y <= pAddPort_1_s_delay_28_Y;
    pAddPort_1_s_delay_29_Z <= pAddPort_1_s_delay_28_Z;
    pAddPort_1_s_delay_29_T <= pAddPort_1_s_delay_28_T;
    pAddPort_1_s_delay_30_X <= pAddPort_1_s_delay_29_X;
    pAddPort_1_s_delay_30_Y <= pAddPort_1_s_delay_29_Y;
    pAddPort_1_s_delay_30_Z <= pAddPort_1_s_delay_29_Z;
    pAddPort_1_s_delay_30_T <= pAddPort_1_s_delay_29_T;
    shiftRegs_addressOutFull_1_delay_1 <= shiftRegs_addressOutFull_1;
    shiftRegs_addressOutFull_1_delay_2 <= shiftRegs_addressOutFull_1_delay_1;
    shiftRegs_addressOutFull_1_delay_3 <= shiftRegs_addressOutFull_1_delay_2;
    shiftRegs_addressOutFull_1_delay_4 <= shiftRegs_addressOutFull_1_delay_3;
    shiftRegs_addressOutFull_1_delay_5 <= shiftRegs_addressOutFull_1_delay_4;
    shiftRegs_addressOutFull_1_delay_6 <= shiftRegs_addressOutFull_1_delay_5;
    shiftRegs_addressOutFull_1_delay_7 <= shiftRegs_addressOutFull_1_delay_6;
    shiftRegs_addressOutFull_1_delay_8 <= shiftRegs_addressOutFull_1_delay_7;
    shiftRegs_addressOutFull_1_delay_9 <= shiftRegs_addressOutFull_1_delay_8;
    shiftRegs_addressOutFull_1_delay_10 <= shiftRegs_addressOutFull_1_delay_9;
    shiftRegs_addressOutFull_1_delay_11 <= shiftRegs_addressOutFull_1_delay_10;
    shiftRegs_addressOutFull_1_delay_12 <= shiftRegs_addressOutFull_1_delay_11;
    shiftRegs_addressOutFull_1_delay_13 <= shiftRegs_addressOutFull_1_delay_12;
    shiftRegs_addressOutFull_1_delay_14 <= shiftRegs_addressOutFull_1_delay_13;
    shiftRegs_addressOutFull_1_delay_15 <= shiftRegs_addressOutFull_1_delay_14;
    shiftRegs_addressOutFull_1_delay_16 <= shiftRegs_addressOutFull_1_delay_15;
    shiftRegs_addressOutFull_1_delay_17 <= shiftRegs_addressOutFull_1_delay_16;
    shiftRegs_addressOutFull_1_delay_18 <= shiftRegs_addressOutFull_1_delay_17;
    shiftRegs_addressOutFull_1_delay_19 <= shiftRegs_addressOutFull_1_delay_18;
    shiftRegs_addressOutFull_1_delay_20 <= shiftRegs_addressOutFull_1_delay_19;
    shiftRegs_addressOutFull_1_delay_21 <= shiftRegs_addressOutFull_1_delay_20;
    shiftRegs_addressOutFull_1_delay_22 <= shiftRegs_addressOutFull_1_delay_21;
    shiftRegs_addressOutFull_1_delay_23 <= shiftRegs_addressOutFull_1_delay_22;
    shiftRegs_addressOutFull_1_delay_24 <= shiftRegs_addressOutFull_1_delay_23;
    shiftRegs_addressOutFull_1_delay_25 <= shiftRegs_addressOutFull_1_delay_24;
    shiftRegs_addressOutFull_1_delay_26 <= shiftRegs_addressOutFull_1_delay_25;
    shiftRegs_addressOutFull_1_delay_27 <= shiftRegs_addressOutFull_1_delay_26;
    shiftRegs_addressOutFull_1_delay_28 <= shiftRegs_addressOutFull_1_delay_27;
    shiftRegs_addressOutFull_1_delay_29 <= shiftRegs_addressOutFull_1_delay_28;
    shiftRegs_addressOutFull_1_delay_30 <= shiftRegs_addressOutFull_1_delay_29;
    stage1_inputData_1_delay_1_X_2 <= stage1_inputData_1_X;
    stage1_inputData_1_delay_1_Y_2 <= stage1_inputData_1_Y;
    stage1_inputData_1_delay_1_Z_2 <= stage1_inputData_1_Z;
    stage1_inputData_1_delay_1_T_2 <= stage1_inputData_1_T;
    stage1_inputData_1_delay_2_X_2 <= stage1_inputData_1_delay_1_X_2;
    stage1_inputData_1_delay_2_Y_2 <= stage1_inputData_1_delay_1_Y_2;
    stage1_inputData_1_delay_2_Z_2 <= stage1_inputData_1_delay_1_Z_2;
    stage1_inputData_1_delay_2_T_2 <= stage1_inputData_1_delay_1_T_2;
    stage1_inputData_1_delay_3_X_2 <= stage1_inputData_1_delay_2_X_2;
    stage1_inputData_1_delay_3_Y_2 <= stage1_inputData_1_delay_2_Y_2;
    stage1_inputData_1_delay_3_Z_2 <= stage1_inputData_1_delay_2_Z_2;
    stage1_inputData_1_delay_3_T_2 <= stage1_inputData_1_delay_2_T_2;
    stage1_inputData_1_delay_4_X_2 <= stage1_inputData_1_delay_3_X_2;
    stage1_inputData_1_delay_4_Y_2 <= stage1_inputData_1_delay_3_Y_2;
    stage1_inputData_1_delay_4_Z_2 <= stage1_inputData_1_delay_3_Z_2;
    stage1_inputData_1_delay_4_T_2 <= stage1_inputData_1_delay_3_T_2;
    stage1_inputData_1_delay_5_X_2 <= stage1_inputData_1_delay_4_X_2;
    stage1_inputData_1_delay_5_Y_2 <= stage1_inputData_1_delay_4_Y_2;
    stage1_inputData_1_delay_5_Z_2 <= stage1_inputData_1_delay_4_Z_2;
    stage1_inputData_1_delay_5_T_2 <= stage1_inputData_1_delay_4_T_2;
    stage1_inputData_1_delay_6_X_1 <= stage1_inputData_1_delay_5_X_2;
    stage1_inputData_1_delay_6_Y_1 <= stage1_inputData_1_delay_5_Y_2;
    stage1_inputData_1_delay_6_Z_1 <= stage1_inputData_1_delay_5_Z_2;
    stage1_inputData_1_delay_6_T_1 <= stage1_inputData_1_delay_5_T_2;
    stage1_inputData_1_delay_7_X_1 <= stage1_inputData_1_delay_6_X_1;
    stage1_inputData_1_delay_7_Y_1 <= stage1_inputData_1_delay_6_Y_1;
    stage1_inputData_1_delay_7_Z_1 <= stage1_inputData_1_delay_6_Z_1;
    stage1_inputData_1_delay_7_T_1 <= stage1_inputData_1_delay_6_T_1;
    stage1_inputData_1_delay_8_X_1 <= stage1_inputData_1_delay_7_X_1;
    stage1_inputData_1_delay_8_Y_1 <= stage1_inputData_1_delay_7_Y_1;
    stage1_inputData_1_delay_8_Z_1 <= stage1_inputData_1_delay_7_Z_1;
    stage1_inputData_1_delay_8_T_1 <= stage1_inputData_1_delay_7_T_1;
    stage1_inputData_1_delay_9_X_1 <= stage1_inputData_1_delay_8_X_1;
    stage1_inputData_1_delay_9_Y_1 <= stage1_inputData_1_delay_8_Y_1;
    stage1_inputData_1_delay_9_Z_1 <= stage1_inputData_1_delay_8_Z_1;
    stage1_inputData_1_delay_9_T_1 <= stage1_inputData_1_delay_8_T_1;
    stage1_inputData_1_delay_10_X_1 <= stage1_inputData_1_delay_9_X_1;
    stage1_inputData_1_delay_10_Y_1 <= stage1_inputData_1_delay_9_Y_1;
    stage1_inputData_1_delay_10_Z_1 <= stage1_inputData_1_delay_9_Z_1;
    stage1_inputData_1_delay_10_T_1 <= stage1_inputData_1_delay_9_T_1;
    stage1_inputData_1_delay_11_X_1 <= stage1_inputData_1_delay_10_X_1;
    stage1_inputData_1_delay_11_Y_1 <= stage1_inputData_1_delay_10_Y_1;
    stage1_inputData_1_delay_11_Z_1 <= stage1_inputData_1_delay_10_Z_1;
    stage1_inputData_1_delay_11_T_1 <= stage1_inputData_1_delay_10_T_1;
    stage1_inputData_1_delay_12_X_1 <= stage1_inputData_1_delay_11_X_1;
    stage1_inputData_1_delay_12_Y_1 <= stage1_inputData_1_delay_11_Y_1;
    stage1_inputData_1_delay_12_Z_1 <= stage1_inputData_1_delay_11_Z_1;
    stage1_inputData_1_delay_12_T_1 <= stage1_inputData_1_delay_11_T_1;
    stage1_inputData_1_delay_13_X_1 <= stage1_inputData_1_delay_12_X_1;
    stage1_inputData_1_delay_13_Y_1 <= stage1_inputData_1_delay_12_Y_1;
    stage1_inputData_1_delay_13_Z_1 <= stage1_inputData_1_delay_12_Z_1;
    stage1_inputData_1_delay_13_T_1 <= stage1_inputData_1_delay_12_T_1;
    stage1_inputData_1_delay_14_X_1 <= stage1_inputData_1_delay_13_X_1;
    stage1_inputData_1_delay_14_Y_1 <= stage1_inputData_1_delay_13_Y_1;
    stage1_inputData_1_delay_14_Z_1 <= stage1_inputData_1_delay_13_Z_1;
    stage1_inputData_1_delay_14_T_1 <= stage1_inputData_1_delay_13_T_1;
    stage1_inputData_1_delay_15_X_1 <= stage1_inputData_1_delay_14_X_1;
    stage1_inputData_1_delay_15_Y_1 <= stage1_inputData_1_delay_14_Y_1;
    stage1_inputData_1_delay_15_Z_1 <= stage1_inputData_1_delay_14_Z_1;
    stage1_inputData_1_delay_15_T_1 <= stage1_inputData_1_delay_14_T_1;
    stage1_inputData_1_delay_16_X_1 <= stage1_inputData_1_delay_15_X_1;
    stage1_inputData_1_delay_16_Y_1 <= stage1_inputData_1_delay_15_Y_1;
    stage1_inputData_1_delay_16_Z_1 <= stage1_inputData_1_delay_15_Z_1;
    stage1_inputData_1_delay_16_T_1 <= stage1_inputData_1_delay_15_T_1;
    stage1_inputData_1_delay_17_X_1 <= stage1_inputData_1_delay_16_X_1;
    stage1_inputData_1_delay_17_Y_1 <= stage1_inputData_1_delay_16_Y_1;
    stage1_inputData_1_delay_17_Z_1 <= stage1_inputData_1_delay_16_Z_1;
    stage1_inputData_1_delay_17_T_1 <= stage1_inputData_1_delay_16_T_1;
    stage1_inputData_1_delay_18_X_1 <= stage1_inputData_1_delay_17_X_1;
    stage1_inputData_1_delay_18_Y_1 <= stage1_inputData_1_delay_17_Y_1;
    stage1_inputData_1_delay_18_Z_1 <= stage1_inputData_1_delay_17_Z_1;
    stage1_inputData_1_delay_18_T_1 <= stage1_inputData_1_delay_17_T_1;
    stage1_inputData_1_delay_19_X_1 <= stage1_inputData_1_delay_18_X_1;
    stage1_inputData_1_delay_19_Y_1 <= stage1_inputData_1_delay_18_Y_1;
    stage1_inputData_1_delay_19_Z_1 <= stage1_inputData_1_delay_18_Z_1;
    stage1_inputData_1_delay_19_T_1 <= stage1_inputData_1_delay_18_T_1;
    stage1_inputData_1_delay_20_X_1 <= stage1_inputData_1_delay_19_X_1;
    stage1_inputData_1_delay_20_Y_1 <= stage1_inputData_1_delay_19_Y_1;
    stage1_inputData_1_delay_20_Z_1 <= stage1_inputData_1_delay_19_Z_1;
    stage1_inputData_1_delay_20_T_1 <= stage1_inputData_1_delay_19_T_1;
    stage1_inputData_1_delay_21_X_1 <= stage1_inputData_1_delay_20_X_1;
    stage1_inputData_1_delay_21_Y_1 <= stage1_inputData_1_delay_20_Y_1;
    stage1_inputData_1_delay_21_Z_1 <= stage1_inputData_1_delay_20_Z_1;
    stage1_inputData_1_delay_21_T_1 <= stage1_inputData_1_delay_20_T_1;
    stage1_inputData_1_delay_22_X_1 <= stage1_inputData_1_delay_21_X_1;
    stage1_inputData_1_delay_22_Y_1 <= stage1_inputData_1_delay_21_Y_1;
    stage1_inputData_1_delay_22_Z_1 <= stage1_inputData_1_delay_21_Z_1;
    stage1_inputData_1_delay_22_T_1 <= stage1_inputData_1_delay_21_T_1;
    stage1_inputData_1_delay_23_X_1 <= stage1_inputData_1_delay_22_X_1;
    stage1_inputData_1_delay_23_Y_1 <= stage1_inputData_1_delay_22_Y_1;
    stage1_inputData_1_delay_23_Z_1 <= stage1_inputData_1_delay_22_Z_1;
    stage1_inputData_1_delay_23_T_1 <= stage1_inputData_1_delay_22_T_1;
    stage1_inputData_1_delay_24_X_1 <= stage1_inputData_1_delay_23_X_1;
    stage1_inputData_1_delay_24_Y_1 <= stage1_inputData_1_delay_23_Y_1;
    stage1_inputData_1_delay_24_Z_1 <= stage1_inputData_1_delay_23_Z_1;
    stage1_inputData_1_delay_24_T_1 <= stage1_inputData_1_delay_23_T_1;
    stage1_inputData_1_delay_25_X_1 <= stage1_inputData_1_delay_24_X_1;
    stage1_inputData_1_delay_25_Y_1 <= stage1_inputData_1_delay_24_Y_1;
    stage1_inputData_1_delay_25_Z_1 <= stage1_inputData_1_delay_24_Z_1;
    stage1_inputData_1_delay_25_T_1 <= stage1_inputData_1_delay_24_T_1;
    stage1_inputData_1_delay_26_X_1 <= stage1_inputData_1_delay_25_X_1;
    stage1_inputData_1_delay_26_Y_1 <= stage1_inputData_1_delay_25_Y_1;
    stage1_inputData_1_delay_26_Z_1 <= stage1_inputData_1_delay_25_Z_1;
    stage1_inputData_1_delay_26_T_1 <= stage1_inputData_1_delay_25_T_1;
    stage1_inputData_1_delay_27_X_1 <= stage1_inputData_1_delay_26_X_1;
    stage1_inputData_1_delay_27_Y_1 <= stage1_inputData_1_delay_26_Y_1;
    stage1_inputData_1_delay_27_Z_1 <= stage1_inputData_1_delay_26_Z_1;
    stage1_inputData_1_delay_27_T_1 <= stage1_inputData_1_delay_26_T_1;
    stage1_inputData_1_delay_28_X_1 <= stage1_inputData_1_delay_27_X_1;
    stage1_inputData_1_delay_28_Y_1 <= stage1_inputData_1_delay_27_Y_1;
    stage1_inputData_1_delay_28_Z_1 <= stage1_inputData_1_delay_27_Z_1;
    stage1_inputData_1_delay_28_T_1 <= stage1_inputData_1_delay_27_T_1;
    stage1_inputData_1_delay_29_X_1 <= stage1_inputData_1_delay_28_X_1;
    stage1_inputData_1_delay_29_Y_1 <= stage1_inputData_1_delay_28_Y_1;
    stage1_inputData_1_delay_29_Z_1 <= stage1_inputData_1_delay_28_Z_1;
    stage1_inputData_1_delay_29_T_1 <= stage1_inputData_1_delay_28_T_1;
    stage1_inputData_1_delay_30_X_1 <= stage1_inputData_1_delay_29_X_1;
    stage1_inputData_1_delay_30_Y_1 <= stage1_inputData_1_delay_29_Y_1;
    stage1_inputData_1_delay_30_Z_1 <= stage1_inputData_1_delay_29_Z_1;
    stage1_inputData_1_delay_30_T_1 <= stage1_inputData_1_delay_29_T_1;
    stage1_inputData_1_delay_31_X_1 <= stage1_inputData_1_delay_30_X_1;
    stage1_inputData_1_delay_31_Y_1 <= stage1_inputData_1_delay_30_Y_1;
    stage1_inputData_1_delay_31_Z_1 <= stage1_inputData_1_delay_30_Z_1;
    stage1_inputData_1_delay_31_T_1 <= stage1_inputData_1_delay_30_T_1;
    stage1_inputData_1_delay_32_X_1 <= stage1_inputData_1_delay_31_X_1;
    stage1_inputData_1_delay_32_Y_1 <= stage1_inputData_1_delay_31_Y_1;
    stage1_inputData_1_delay_32_Z_1 <= stage1_inputData_1_delay_31_Z_1;
    stage1_inputData_1_delay_32_T_1 <= stage1_inputData_1_delay_31_T_1;
    stage1_inputData_1_delay_33_X_1 <= stage1_inputData_1_delay_32_X_1;
    stage1_inputData_1_delay_33_Y_1 <= stage1_inputData_1_delay_32_Y_1;
    stage1_inputData_1_delay_33_Z_1 <= stage1_inputData_1_delay_32_Z_1;
    stage1_inputData_1_delay_33_T_1 <= stage1_inputData_1_delay_32_T_1;
    stage1_inputData_1_delay_34_X_1 <= stage1_inputData_1_delay_33_X_1;
    stage1_inputData_1_delay_34_Y_1 <= stage1_inputData_1_delay_33_Y_1;
    stage1_inputData_1_delay_34_Z_1 <= stage1_inputData_1_delay_33_Z_1;
    stage1_inputData_1_delay_34_T_1 <= stage1_inputData_1_delay_33_T_1;
    stage1_inputData_1_delay_35_X_1 <= stage1_inputData_1_delay_34_X_1;
    stage1_inputData_1_delay_35_Y_1 <= stage1_inputData_1_delay_34_Y_1;
    stage1_inputData_1_delay_35_Z_1 <= stage1_inputData_1_delay_34_Z_1;
    stage1_inputData_1_delay_35_T_1 <= stage1_inputData_1_delay_34_T_1;
    stage1_inputAddress_1_delay_1_1 <= stage1_inputAddress_1;
    stage1_inputAddress_1_delay_2_1 <= stage1_inputAddress_1_delay_1_1;
    stage1_inputAddress_1_delay_3_1 <= stage1_inputAddress_1_delay_2_1;
    stage1_inputAddress_1_delay_4_1 <= stage1_inputAddress_1_delay_3_1;
    stage1_inputAddress_1_delay_5_1 <= stage1_inputAddress_1_delay_4_1;
    stage1_inputAddress_1_delay_6 <= stage1_inputAddress_1_delay_5_1;
    stage1_inputAddress_1_delay_7 <= stage1_inputAddress_1_delay_6;
    stage1_inputAddress_1_delay_8 <= stage1_inputAddress_1_delay_7;
    stage1_inputAddress_1_delay_9 <= stage1_inputAddress_1_delay_8;
    stage1_inputAddress_1_delay_10 <= stage1_inputAddress_1_delay_9;
    stage1_inputAddress_1_delay_11 <= stage1_inputAddress_1_delay_10;
    stage1_inputAddress_1_delay_12 <= stage1_inputAddress_1_delay_11;
    stage1_inputAddress_1_delay_13 <= stage1_inputAddress_1_delay_12;
    stage1_inputAddress_1_delay_14 <= stage1_inputAddress_1_delay_13;
    stage1_inputAddress_1_delay_15 <= stage1_inputAddress_1_delay_14;
    stage1_inputAddress_1_delay_16 <= stage1_inputAddress_1_delay_15;
    stage1_inputAddress_1_delay_17 <= stage1_inputAddress_1_delay_16;
    stage1_inputAddress_1_delay_18 <= stage1_inputAddress_1_delay_17;
    stage1_inputAddress_1_delay_19 <= stage1_inputAddress_1_delay_18;
    stage1_inputAddress_1_delay_20 <= stage1_inputAddress_1_delay_19;
    stage1_inputAddress_1_delay_21 <= stage1_inputAddress_1_delay_20;
    stage1_inputAddress_1_delay_22 <= stage1_inputAddress_1_delay_21;
    stage1_inputAddress_1_delay_23 <= stage1_inputAddress_1_delay_22;
    stage1_inputAddress_1_delay_24 <= stage1_inputAddress_1_delay_23;
    stage1_inputAddress_1_delay_25 <= stage1_inputAddress_1_delay_24;
    stage1_inputAddress_1_delay_26 <= stage1_inputAddress_1_delay_25;
    stage1_inputAddress_1_delay_27 <= stage1_inputAddress_1_delay_26;
    stage1_inputAddress_1_delay_28 <= stage1_inputAddress_1_delay_27;
    stage1_inputAddress_1_delay_29 <= stage1_inputAddress_1_delay_28;
    stage1_inputAddress_1_delay_30 <= stage1_inputAddress_1_delay_29;
    stage1_inputAddress_1_delay_31 <= stage1_inputAddress_1_delay_30;
    stage1_inputAddress_1_delay_32 <= stage1_inputAddress_1_delay_31;
    stage1_inputAddress_1_delay_33 <= stage1_inputAddress_1_delay_32;
    stage1_inputAddress_1_delay_34 <= stage1_inputAddress_1_delay_33;
    stage1_inputAddress_1_delay_35 <= stage1_inputAddress_1_delay_34;
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      _zz_io_dataIn_0_valid_5 <= 1'b0;
      _zz_io_dataIn_0_valid_6 <= 1'b0;
      _zz_io_dataIn_0_valid_7 <= 1'b0;
      _zz_io_dataIn_0_valid_8 <= 1'b0;
      _zz_io_dataIn_0_valid_9 <= 1'b0;
      _zz_io_dataIn_0_valid_10 <= 1'b0;
      _zz_io_dataIn_0_valid_11 <= 1'b0;
      _zz_io_dataIn_0_valid_12 <= 1'b0;
      _zz_io_dataIn_0_valid_13 <= 1'b0;
      _zz_io_dataIn_0_valid_14 <= 1'b0;
      _zz_io_dataIn_0_valid_15 <= 1'b0;
      _zz_io_dataIn_0_valid_16 <= 1'b0;
      _zz_io_dataIn_0_valid_17 <= 1'b0;
      _zz_io_dataIn_0_valid_18 <= 1'b0;
      _zz_io_dataIn_0_valid_19 <= 1'b0;
      _zz_io_dataIn_0_valid_20 <= 1'b0;
      _zz_io_dataIn_0_valid_21 <= 1'b0;
      _zz_io_dataIn_0_valid_22 <= 1'b0;
      _zz_io_dataIn_0_valid_23 <= 1'b0;
      _zz_io_dataIn_0_valid_24 <= 1'b0;
      _zz_io_dataIn_0_valid_25 <= 1'b0;
      _zz_io_dataIn_0_valid_26 <= 1'b0;
      _zz_io_dataIn_0_valid_27 <= 1'b0;
      _zz_io_dataIn_0_valid_28 <= 1'b0;
      _zz_io_dataIn_0_valid_29 <= 1'b0;
      _zz_io_dataIn_0_valid_30 <= 1'b0;
      _zz_io_dataIn_0_valid_31 <= 1'b0;
      _zz_io_dataIn_0_valid_32 <= 1'b0;
      _zz_io_dataIn_0_valid_33 <= 1'b0;
      _zz_io_dataIn_0_valid_34 <= 1'b0;
      _zz_io_dataIn_1_valid <= 1'b0;
      _zz_io_dataIn_1_valid_1 <= 1'b0;
      _zz_io_dataIn_1_valid_2 <= 1'b0;
      _zz_io_dataIn_1_valid_3 <= 1'b0;
      _zz_io_dataIn_1_valid_4 <= 1'b0;
      _zz_io_dataIn_1_valid_5 <= 1'b0;
      _zz_io_dataIn_1_valid_6 <= 1'b0;
      _zz_io_dataIn_1_valid_7 <= 1'b0;
      _zz_io_dataIn_1_valid_8 <= 1'b0;
      _zz_io_dataIn_1_valid_9 <= 1'b0;
      _zz_io_dataIn_1_valid_10 <= 1'b0;
      _zz_io_dataIn_1_valid_11 <= 1'b0;
      _zz_io_dataIn_1_valid_12 <= 1'b0;
      _zz_io_dataIn_1_valid_13 <= 1'b0;
      _zz_io_dataIn_1_valid_14 <= 1'b0;
      _zz_io_dataIn_1_valid_15 <= 1'b0;
      _zz_io_dataIn_1_valid_16 <= 1'b0;
      _zz_io_dataIn_1_valid_17 <= 1'b0;
      _zz_io_dataIn_1_valid_18 <= 1'b0;
      _zz_io_dataIn_1_valid_19 <= 1'b0;
      _zz_io_dataIn_1_valid_20 <= 1'b0;
      _zz_io_dataIn_1_valid_21 <= 1'b0;
      _zz_io_dataIn_1_valid_22 <= 1'b0;
      _zz_io_dataIn_1_valid_23 <= 1'b0;
      _zz_io_dataIn_1_valid_24 <= 1'b0;
      _zz_io_dataIn_1_valid_25 <= 1'b0;
      _zz_io_dataIn_1_valid_26 <= 1'b0;
      _zz_io_dataIn_1_valid_27 <= 1'b0;
      _zz_io_dataIn_1_valid_28 <= 1'b0;
      _zz_io_dataIn_1_valid_29 <= 1'b0;
      _zz_io_dataIn_1_valid_30 <= 1'b0;
      _zz_io_dataIn_1_valid_31 <= 1'b0;
      _zz_io_dataIn_1_valid_32 <= 1'b0;
      _zz_io_dataIn_1_valid_33 <= 1'b0;
      _zz_io_dataIn_1_valid_34 <= 1'b0;
      _zz_io_dataIn_0_valid_40 <= 1'b0;
      _zz_io_dataIn_0_valid_41 <= 1'b0;
      _zz_io_dataIn_0_valid_42 <= 1'b0;
      _zz_io_dataIn_0_valid_43 <= 1'b0;
      _zz_io_dataIn_0_valid_44 <= 1'b0;
      _zz_io_dataIn_0_valid_45 <= 1'b0;
      _zz_io_dataIn_0_valid_46 <= 1'b0;
      _zz_io_dataIn_0_valid_47 <= 1'b0;
      _zz_io_dataIn_0_valid_48 <= 1'b0;
      _zz_io_dataIn_0_valid_49 <= 1'b0;
      _zz_io_dataIn_0_valid_50 <= 1'b0;
      _zz_io_dataIn_0_valid_51 <= 1'b0;
      _zz_io_dataIn_0_valid_52 <= 1'b0;
      _zz_io_dataIn_0_valid_53 <= 1'b0;
      _zz_io_dataIn_0_valid_54 <= 1'b0;
      _zz_io_dataIn_0_valid_55 <= 1'b0;
      _zz_io_dataIn_0_valid_56 <= 1'b0;
      _zz_io_dataIn_0_valid_57 <= 1'b0;
      _zz_io_dataIn_0_valid_58 <= 1'b0;
      _zz_io_dataIn_0_valid_59 <= 1'b0;
      _zz_io_dataIn_0_valid_60 <= 1'b0;
      _zz_io_dataIn_0_valid_61 <= 1'b0;
      _zz_io_dataIn_0_valid_62 <= 1'b0;
      _zz_io_dataIn_0_valid_63 <= 1'b0;
      _zz_io_dataIn_0_valid_64 <= 1'b0;
      _zz_io_dataIn_0_valid_65 <= 1'b0;
      _zz_io_dataIn_0_valid_66 <= 1'b0;
      _zz_io_dataIn_0_valid_67 <= 1'b0;
      _zz_io_dataIn_0_valid_68 <= 1'b0;
      _zz_io_dataIn_0_valid_69 <= 1'b0;
      _zz_io_dataIn_1_valid_35 <= 1'b0;
      _zz_io_dataIn_1_valid_36 <= 1'b0;
      _zz_io_dataIn_1_valid_37 <= 1'b0;
      _zz_io_dataIn_1_valid_38 <= 1'b0;
      _zz_io_dataIn_1_valid_39 <= 1'b0;
      _zz_io_dataIn_1_valid_40 <= 1'b0;
      _zz_io_dataIn_1_valid_41 <= 1'b0;
      _zz_io_dataIn_1_valid_42 <= 1'b0;
      _zz_io_dataIn_1_valid_43 <= 1'b0;
      _zz_io_dataIn_1_valid_44 <= 1'b0;
      _zz_io_dataIn_1_valid_45 <= 1'b0;
      _zz_io_dataIn_1_valid_46 <= 1'b0;
      _zz_io_dataIn_1_valid_47 <= 1'b0;
      _zz_io_dataIn_1_valid_48 <= 1'b0;
      _zz_io_dataIn_1_valid_49 <= 1'b0;
      _zz_io_dataIn_1_valid_50 <= 1'b0;
      _zz_io_dataIn_1_valid_51 <= 1'b0;
      _zz_io_dataIn_1_valid_52 <= 1'b0;
      _zz_io_dataIn_1_valid_53 <= 1'b0;
      _zz_io_dataIn_1_valid_54 <= 1'b0;
      _zz_io_dataIn_1_valid_55 <= 1'b0;
      _zz_io_dataIn_1_valid_56 <= 1'b0;
      _zz_io_dataIn_1_valid_57 <= 1'b0;
      _zz_io_dataIn_1_valid_58 <= 1'b0;
      _zz_io_dataIn_1_valid_59 <= 1'b0;
      _zz_io_dataIn_1_valid_60 <= 1'b0;
      _zz_io_dataIn_1_valid_61 <= 1'b0;
      _zz_io_dataIn_1_valid_62 <= 1'b0;
      _zz_io_dataIn_1_valid_63 <= 1'b0;
      _zz_io_dataIn_1_valid_64 <= 1'b0;
      _zz_io_dataIn_1_valid_65 <= 1'b0;
      _zz_io_dataIn_1_valid_66 <= 1'b0;
      _zz_io_dataIn_1_valid_67 <= 1'b0;
      _zz_io_dataIn_1_valid_68 <= 1'b0;
      _zz_io_dataIn_1_valid_69 <= 1'b0;
    end else begin
      _zz_io_dataIn_0_valid_5 <= ((stateRam_0_io_state_0 || _zz_io_dataIn_0_valid_4) && shiftRegs_validOutFull_0);
      _zz_io_dataIn_0_valid_6 <= _zz_io_dataIn_0_valid_5;
      _zz_io_dataIn_0_valid_7 <= _zz_io_dataIn_0_valid_6;
      _zz_io_dataIn_0_valid_8 <= _zz_io_dataIn_0_valid_7;
      _zz_io_dataIn_0_valid_9 <= _zz_io_dataIn_0_valid_8;
      _zz_io_dataIn_0_valid_10 <= _zz_io_dataIn_0_valid_9;
      _zz_io_dataIn_0_valid_11 <= _zz_io_dataIn_0_valid_10;
      _zz_io_dataIn_0_valid_12 <= _zz_io_dataIn_0_valid_11;
      _zz_io_dataIn_0_valid_13 <= _zz_io_dataIn_0_valid_12;
      _zz_io_dataIn_0_valid_14 <= _zz_io_dataIn_0_valid_13;
      _zz_io_dataIn_0_valid_15 <= _zz_io_dataIn_0_valid_14;
      _zz_io_dataIn_0_valid_16 <= _zz_io_dataIn_0_valid_15;
      _zz_io_dataIn_0_valid_17 <= _zz_io_dataIn_0_valid_16;
      _zz_io_dataIn_0_valid_18 <= _zz_io_dataIn_0_valid_17;
      _zz_io_dataIn_0_valid_19 <= _zz_io_dataIn_0_valid_18;
      _zz_io_dataIn_0_valid_20 <= _zz_io_dataIn_0_valid_19;
      _zz_io_dataIn_0_valid_21 <= _zz_io_dataIn_0_valid_20;
      _zz_io_dataIn_0_valid_22 <= _zz_io_dataIn_0_valid_21;
      _zz_io_dataIn_0_valid_23 <= _zz_io_dataIn_0_valid_22;
      _zz_io_dataIn_0_valid_24 <= _zz_io_dataIn_0_valid_23;
      _zz_io_dataIn_0_valid_25 <= _zz_io_dataIn_0_valid_24;
      _zz_io_dataIn_0_valid_26 <= _zz_io_dataIn_0_valid_25;
      _zz_io_dataIn_0_valid_27 <= _zz_io_dataIn_0_valid_26;
      _zz_io_dataIn_0_valid_28 <= _zz_io_dataIn_0_valid_27;
      _zz_io_dataIn_0_valid_29 <= _zz_io_dataIn_0_valid_28;
      _zz_io_dataIn_0_valid_30 <= _zz_io_dataIn_0_valid_29;
      _zz_io_dataIn_0_valid_31 <= _zz_io_dataIn_0_valid_30;
      _zz_io_dataIn_0_valid_32 <= _zz_io_dataIn_0_valid_31;
      _zz_io_dataIn_0_valid_33 <= _zz_io_dataIn_0_valid_32;
      _zz_io_dataIn_0_valid_34 <= _zz_io_dataIn_0_valid_33;
      _zz_io_dataIn_1_valid <= (stage1_inputValid_0 && (! (shiftRegs_validOut_0 && (stage1_inputAddress_0 == shiftRegs_addressOut_0))));
      _zz_io_dataIn_1_valid_1 <= _zz_io_dataIn_1_valid;
      _zz_io_dataIn_1_valid_2 <= _zz_io_dataIn_1_valid_1;
      _zz_io_dataIn_1_valid_3 <= _zz_io_dataIn_1_valid_2;
      _zz_io_dataIn_1_valid_4 <= _zz_io_dataIn_1_valid_3;
      _zz_io_dataIn_1_valid_5 <= (stateRam_0_io_state_1 && _zz_io_dataIn_1_valid_4);
      _zz_io_dataIn_1_valid_6 <= _zz_io_dataIn_1_valid_5;
      _zz_io_dataIn_1_valid_7 <= _zz_io_dataIn_1_valid_6;
      _zz_io_dataIn_1_valid_8 <= _zz_io_dataIn_1_valid_7;
      _zz_io_dataIn_1_valid_9 <= _zz_io_dataIn_1_valid_8;
      _zz_io_dataIn_1_valid_10 <= _zz_io_dataIn_1_valid_9;
      _zz_io_dataIn_1_valid_11 <= _zz_io_dataIn_1_valid_10;
      _zz_io_dataIn_1_valid_12 <= _zz_io_dataIn_1_valid_11;
      _zz_io_dataIn_1_valid_13 <= _zz_io_dataIn_1_valid_12;
      _zz_io_dataIn_1_valid_14 <= _zz_io_dataIn_1_valid_13;
      _zz_io_dataIn_1_valid_15 <= _zz_io_dataIn_1_valid_14;
      _zz_io_dataIn_1_valid_16 <= _zz_io_dataIn_1_valid_15;
      _zz_io_dataIn_1_valid_17 <= _zz_io_dataIn_1_valid_16;
      _zz_io_dataIn_1_valid_18 <= _zz_io_dataIn_1_valid_17;
      _zz_io_dataIn_1_valid_19 <= _zz_io_dataIn_1_valid_18;
      _zz_io_dataIn_1_valid_20 <= _zz_io_dataIn_1_valid_19;
      _zz_io_dataIn_1_valid_21 <= _zz_io_dataIn_1_valid_20;
      _zz_io_dataIn_1_valid_22 <= _zz_io_dataIn_1_valid_21;
      _zz_io_dataIn_1_valid_23 <= _zz_io_dataIn_1_valid_22;
      _zz_io_dataIn_1_valid_24 <= _zz_io_dataIn_1_valid_23;
      _zz_io_dataIn_1_valid_25 <= _zz_io_dataIn_1_valid_24;
      _zz_io_dataIn_1_valid_26 <= _zz_io_dataIn_1_valid_25;
      _zz_io_dataIn_1_valid_27 <= _zz_io_dataIn_1_valid_26;
      _zz_io_dataIn_1_valid_28 <= _zz_io_dataIn_1_valid_27;
      _zz_io_dataIn_1_valid_29 <= _zz_io_dataIn_1_valid_28;
      _zz_io_dataIn_1_valid_30 <= _zz_io_dataIn_1_valid_29;
      _zz_io_dataIn_1_valid_31 <= _zz_io_dataIn_1_valid_30;
      _zz_io_dataIn_1_valid_32 <= _zz_io_dataIn_1_valid_31;
      _zz_io_dataIn_1_valid_33 <= _zz_io_dataIn_1_valid_32;
      _zz_io_dataIn_1_valid_34 <= _zz_io_dataIn_1_valid_33;
      _zz_io_dataIn_0_valid_40 <= ((stateRam_1_1_io_state_0 || _zz_io_dataIn_0_valid_39) && shiftRegs_validOutFull_1);
      _zz_io_dataIn_0_valid_41 <= _zz_io_dataIn_0_valid_40;
      _zz_io_dataIn_0_valid_42 <= _zz_io_dataIn_0_valid_41;
      _zz_io_dataIn_0_valid_43 <= _zz_io_dataIn_0_valid_42;
      _zz_io_dataIn_0_valid_44 <= _zz_io_dataIn_0_valid_43;
      _zz_io_dataIn_0_valid_45 <= _zz_io_dataIn_0_valid_44;
      _zz_io_dataIn_0_valid_46 <= _zz_io_dataIn_0_valid_45;
      _zz_io_dataIn_0_valid_47 <= _zz_io_dataIn_0_valid_46;
      _zz_io_dataIn_0_valid_48 <= _zz_io_dataIn_0_valid_47;
      _zz_io_dataIn_0_valid_49 <= _zz_io_dataIn_0_valid_48;
      _zz_io_dataIn_0_valid_50 <= _zz_io_dataIn_0_valid_49;
      _zz_io_dataIn_0_valid_51 <= _zz_io_dataIn_0_valid_50;
      _zz_io_dataIn_0_valid_52 <= _zz_io_dataIn_0_valid_51;
      _zz_io_dataIn_0_valid_53 <= _zz_io_dataIn_0_valid_52;
      _zz_io_dataIn_0_valid_54 <= _zz_io_dataIn_0_valid_53;
      _zz_io_dataIn_0_valid_55 <= _zz_io_dataIn_0_valid_54;
      _zz_io_dataIn_0_valid_56 <= _zz_io_dataIn_0_valid_55;
      _zz_io_dataIn_0_valid_57 <= _zz_io_dataIn_0_valid_56;
      _zz_io_dataIn_0_valid_58 <= _zz_io_dataIn_0_valid_57;
      _zz_io_dataIn_0_valid_59 <= _zz_io_dataIn_0_valid_58;
      _zz_io_dataIn_0_valid_60 <= _zz_io_dataIn_0_valid_59;
      _zz_io_dataIn_0_valid_61 <= _zz_io_dataIn_0_valid_60;
      _zz_io_dataIn_0_valid_62 <= _zz_io_dataIn_0_valid_61;
      _zz_io_dataIn_0_valid_63 <= _zz_io_dataIn_0_valid_62;
      _zz_io_dataIn_0_valid_64 <= _zz_io_dataIn_0_valid_63;
      _zz_io_dataIn_0_valid_65 <= _zz_io_dataIn_0_valid_64;
      _zz_io_dataIn_0_valid_66 <= _zz_io_dataIn_0_valid_65;
      _zz_io_dataIn_0_valid_67 <= _zz_io_dataIn_0_valid_66;
      _zz_io_dataIn_0_valid_68 <= _zz_io_dataIn_0_valid_67;
      _zz_io_dataIn_0_valid_69 <= _zz_io_dataIn_0_valid_68;
      _zz_io_dataIn_1_valid_35 <= (stage1_inputValid_1 && (! (shiftRegs_validOut_1 && (stage1_inputAddress_1 == shiftRegs_addressOut_1))));
      _zz_io_dataIn_1_valid_36 <= _zz_io_dataIn_1_valid_35;
      _zz_io_dataIn_1_valid_37 <= _zz_io_dataIn_1_valid_36;
      _zz_io_dataIn_1_valid_38 <= _zz_io_dataIn_1_valid_37;
      _zz_io_dataIn_1_valid_39 <= _zz_io_dataIn_1_valid_38;
      _zz_io_dataIn_1_valid_40 <= (stateRam_1_1_io_state_1 && _zz_io_dataIn_1_valid_39);
      _zz_io_dataIn_1_valid_41 <= _zz_io_dataIn_1_valid_40;
      _zz_io_dataIn_1_valid_42 <= _zz_io_dataIn_1_valid_41;
      _zz_io_dataIn_1_valid_43 <= _zz_io_dataIn_1_valid_42;
      _zz_io_dataIn_1_valid_44 <= _zz_io_dataIn_1_valid_43;
      _zz_io_dataIn_1_valid_45 <= _zz_io_dataIn_1_valid_44;
      _zz_io_dataIn_1_valid_46 <= _zz_io_dataIn_1_valid_45;
      _zz_io_dataIn_1_valid_47 <= _zz_io_dataIn_1_valid_46;
      _zz_io_dataIn_1_valid_48 <= _zz_io_dataIn_1_valid_47;
      _zz_io_dataIn_1_valid_49 <= _zz_io_dataIn_1_valid_48;
      _zz_io_dataIn_1_valid_50 <= _zz_io_dataIn_1_valid_49;
      _zz_io_dataIn_1_valid_51 <= _zz_io_dataIn_1_valid_50;
      _zz_io_dataIn_1_valid_52 <= _zz_io_dataIn_1_valid_51;
      _zz_io_dataIn_1_valid_53 <= _zz_io_dataIn_1_valid_52;
      _zz_io_dataIn_1_valid_54 <= _zz_io_dataIn_1_valid_53;
      _zz_io_dataIn_1_valid_55 <= _zz_io_dataIn_1_valid_54;
      _zz_io_dataIn_1_valid_56 <= _zz_io_dataIn_1_valid_55;
      _zz_io_dataIn_1_valid_57 <= _zz_io_dataIn_1_valid_56;
      _zz_io_dataIn_1_valid_58 <= _zz_io_dataIn_1_valid_57;
      _zz_io_dataIn_1_valid_59 <= _zz_io_dataIn_1_valid_58;
      _zz_io_dataIn_1_valid_60 <= _zz_io_dataIn_1_valid_59;
      _zz_io_dataIn_1_valid_61 <= _zz_io_dataIn_1_valid_60;
      _zz_io_dataIn_1_valid_62 <= _zz_io_dataIn_1_valid_61;
      _zz_io_dataIn_1_valid_63 <= _zz_io_dataIn_1_valid_62;
      _zz_io_dataIn_1_valid_64 <= _zz_io_dataIn_1_valid_63;
      _zz_io_dataIn_1_valid_65 <= _zz_io_dataIn_1_valid_64;
      _zz_io_dataIn_1_valid_66 <= _zz_io_dataIn_1_valid_65;
      _zz_io_dataIn_1_valid_67 <= _zz_io_dataIn_1_valid_66;
      _zz_io_dataIn_1_valid_68 <= _zz_io_dataIn_1_valid_67;
      _zz_io_dataIn_1_valid_69 <= _zz_io_dataIn_1_valid_68;
    end
  end

  always @(posedge clk) begin
    _zz_io_state_1 <= (stage2_wCnt_value == 12'hfff);
    _zz_io_state_1_1 <= _zz_io_state_1;
    _zz_io_state_1_2 <= _zz_io_state_1_1;
    _zz_io_state_1_3 <= _zz_io_state_1_2;
    _zz_io_state_1_4 <= _zz_io_state_1_3;
    _zz_io_state_1_5 <= (! stage2_calCnt_value[1]);
    _zz_io_state_1_6 <= _zz_io_state_1_5;
    _zz_io_state_1_7 <= _zz_io_state_1_6;
    _zz_io_state_1_8 <= _zz_io_state_1_7;
    _zz_io_state_1_9 <= _zz_io_state_1_8;
    _zz_io_state_1_10 <= (|stage2_calCnt_value);
    _zz_io_state_1_11 <= _zz_io_state_1_10;
    _zz_io_state_1_12 <= _zz_io_state_1_11;
    _zz_io_state_1_13 <= _zz_io_state_1_12;
    _zz_io_state_1_14 <= _zz_io_state_1_13;
    _zz_io_state_1_15 <= (_zz_io_state_1_4 ? (_zz_io_state_1_9 && stateRam_0_io_state_0) : (_zz_io_state_1_14 || stateRam_0_io_state_0));
    _zz_io_state_1_16 <= _zz_io_state_1_15;
    _zz_io_state_1_17 <= _zz_io_state_1_16;
    _zz_io_state_1_18 <= _zz_io_state_1_17;
    _zz_io_state_1_19 <= _zz_io_state_1_18;
    _zz_io_state_1_20 <= _zz_io_state_1_19;
    _zz_io_state_1_21 <= _zz_io_state_1_20;
    _zz_io_state_1_22 <= _zz_io_state_1_21;
    _zz_io_state_1_23 <= _zz_io_state_1_22;
    _zz_io_state_1_24 <= _zz_io_state_1_23;
    _zz_io_state_1_25 <= _zz_io_state_1_24;
    _zz_io_state_1_26 <= _zz_io_state_1_25;
    _zz_io_state_1_27 <= _zz_io_state_1_26;
    _zz_io_state_1_28 <= _zz_io_state_1_27;
    _zz_io_state_1_29 <= _zz_io_state_1_28;
    _zz_io_state_1_30 <= _zz_io_state_1_29;
    _zz_io_state_1_31 <= _zz_io_state_1_30;
    _zz_io_state_1_32 <= _zz_io_state_1_31;
    _zz_io_state_1_33 <= _zz_io_state_1_32;
    _zz_io_state_1_34 <= _zz_io_state_1_33;
    _zz_io_state_1_35 <= _zz_io_state_1_34;
    _zz_io_state_1_36 <= _zz_io_state_1_35;
    _zz_io_state_1_37 <= _zz_io_state_1_36;
    _zz_io_state_1_38 <= _zz_io_state_1_37;
    pippenger_1_dataRam_0_io_rData_1_regNext_X <= dataRam_0_io_rData_1_X;
    pippenger_1_dataRam_0_io_rData_1_regNext_Y <= dataRam_0_io_rData_1_Y;
    pippenger_1_dataRam_0_io_rData_1_regNext_Z <= dataRam_0_io_rData_1_Z;
    pippenger_1_dataRam_0_io_rData_1_regNext_T <= dataRam_0_io_rData_1_T;
    _zz_io_dataIn_1_payload_address <= {stage2_GCnt_value,_zz__zz_io_dataIn_1_payload_address};
    _zz_io_dataIn_1_payload_address_1 <= _zz_io_dataIn_1_payload_address;
    _zz_io_dataIn_1_payload_address_2 <= _zz_io_dataIn_1_payload_address_1;
    _zz_io_dataIn_1_payload_address_3 <= _zz_io_dataIn_1_payload_address_2;
    _zz_io_dataIn_1_payload_address_4 <= _zz_io_dataIn_1_payload_address_3;
    _zz_io_dataIn_1_payload_address_5 <= _zz_io_dataIn_1_payload_address_4;
    _zz_io_dataIn_1_payload_address_6 <= _zz_io_dataIn_1_payload_address_5;
    _zz_io_dataIn_1_payload_address_7 <= _zz_io_dataIn_1_payload_address_6;
    _zz_io_dataIn_1_payload_address_8 <= _zz_io_dataIn_1_payload_address_7;
    _zz_io_dataIn_1_payload_address_9 <= _zz_io_dataIn_1_payload_address_8;
    _zz_io_dataIn_1_payload_address_10 <= _zz_io_dataIn_1_payload_address_9;
    _zz_io_dataIn_1_payload_address_11 <= _zz_io_dataIn_1_payload_address_10;
    _zz_io_dataIn_1_payload_address_12 <= _zz_io_dataIn_1_payload_address_11;
    _zz_io_dataIn_1_payload_address_13 <= _zz_io_dataIn_1_payload_address_12;
    _zz_io_dataIn_1_payload_address_14 <= _zz_io_dataIn_1_payload_address_13;
    _zz_io_dataIn_1_payload_address_15 <= _zz_io_dataIn_1_payload_address_14;
    _zz_io_dataIn_1_payload_address_16 <= _zz_io_dataIn_1_payload_address_15;
    _zz_io_dataIn_1_payload_address_17 <= _zz_io_dataIn_1_payload_address_16;
    _zz_io_dataIn_1_payload_address_18 <= _zz_io_dataIn_1_payload_address_17;
    _zz_io_dataIn_1_payload_address_19 <= _zz_io_dataIn_1_payload_address_18;
    _zz_io_dataIn_1_payload_address_20 <= _zz_io_dataIn_1_payload_address_19;
    _zz_io_dataIn_1_payload_address_21 <= _zz_io_dataIn_1_payload_address_20;
    _zz_io_dataIn_1_payload_address_22 <= _zz_io_dataIn_1_payload_address_21;
    _zz_io_dataIn_1_payload_address_23 <= _zz_io_dataIn_1_payload_address_22;
    _zz_io_dataIn_1_payload_address_24 <= _zz_io_dataIn_1_payload_address_23;
    _zz_io_dataIn_1_payload_address_25 <= _zz_io_dataIn_1_payload_address_24;
    _zz_io_dataIn_1_payload_address_26 <= _zz_io_dataIn_1_payload_address_25;
    _zz_io_dataIn_1_payload_address_27 <= _zz_io_dataIn_1_payload_address_26;
    _zz_io_dataIn_1_payload_address_28 <= _zz_io_dataIn_1_payload_address_27;
    _zz_io_dataIn_1_payload_address_29 <= _zz_io_dataIn_1_payload_address_28;
    _zz_io_state_1_39 <= (stage2_wCnt_value == 12'hfff);
    _zz_io_state_1_40 <= _zz_io_state_1_39;
    _zz_io_state_1_41 <= _zz_io_state_1_40;
    _zz_io_state_1_42 <= _zz_io_state_1_41;
    _zz_io_state_1_43 <= _zz_io_state_1_42;
    _zz_io_state_1_44 <= (! stage2_calCnt_value[1]);
    _zz_io_state_1_45 <= _zz_io_state_1_44;
    _zz_io_state_1_46 <= _zz_io_state_1_45;
    _zz_io_state_1_47 <= _zz_io_state_1_46;
    _zz_io_state_1_48 <= _zz_io_state_1_47;
    _zz_io_state_1_49 <= (|stage2_calCnt_value);
    _zz_io_state_1_50 <= _zz_io_state_1_49;
    _zz_io_state_1_51 <= _zz_io_state_1_50;
    _zz_io_state_1_52 <= _zz_io_state_1_51;
    _zz_io_state_1_53 <= _zz_io_state_1_52;
    _zz_io_state_1_54 <= (_zz_io_state_1_43 ? (_zz_io_state_1_48 && stateRam_1_1_io_state_0) : (_zz_io_state_1_53 || stateRam_1_1_io_state_0));
    _zz_io_state_1_55 <= _zz_io_state_1_54;
    _zz_io_state_1_56 <= _zz_io_state_1_55;
    _zz_io_state_1_57 <= _zz_io_state_1_56;
    _zz_io_state_1_58 <= _zz_io_state_1_57;
    _zz_io_state_1_59 <= _zz_io_state_1_58;
    _zz_io_state_1_60 <= _zz_io_state_1_59;
    _zz_io_state_1_61 <= _zz_io_state_1_60;
    _zz_io_state_1_62 <= _zz_io_state_1_61;
    _zz_io_state_1_63 <= _zz_io_state_1_62;
    _zz_io_state_1_64 <= _zz_io_state_1_63;
    _zz_io_state_1_65 <= _zz_io_state_1_64;
    _zz_io_state_1_66 <= _zz_io_state_1_65;
    _zz_io_state_1_67 <= _zz_io_state_1_66;
    _zz_io_state_1_68 <= _zz_io_state_1_67;
    _zz_io_state_1_69 <= _zz_io_state_1_68;
    _zz_io_state_1_70 <= _zz_io_state_1_69;
    _zz_io_state_1_71 <= _zz_io_state_1_70;
    _zz_io_state_1_72 <= _zz_io_state_1_71;
    _zz_io_state_1_73 <= _zz_io_state_1_72;
    _zz_io_state_1_74 <= _zz_io_state_1_73;
    _zz_io_state_1_75 <= _zz_io_state_1_74;
    _zz_io_state_1_76 <= _zz_io_state_1_75;
    _zz_io_state_1_77 <= _zz_io_state_1_76;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_X <= dataRam_1_1_io_rData_1_X;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_Y <= dataRam_1_1_io_rData_1_Y;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_Z <= dataRam_1_1_io_rData_1_Z;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_T <= dataRam_1_1_io_rData_1_T;
    _zz_io_dataIn_1_payload_address_30 <= {stage2_GCnt_value,_zz__zz_io_dataIn_1_payload_address_30};
    _zz_io_dataIn_1_payload_address_31 <= _zz_io_dataIn_1_payload_address_30;
    _zz_io_dataIn_1_payload_address_32 <= _zz_io_dataIn_1_payload_address_31;
    _zz_io_dataIn_1_payload_address_33 <= _zz_io_dataIn_1_payload_address_32;
    _zz_io_dataIn_1_payload_address_34 <= _zz_io_dataIn_1_payload_address_33;
    _zz_io_dataIn_1_payload_address_35 <= _zz_io_dataIn_1_payload_address_34;
    _zz_io_dataIn_1_payload_address_36 <= _zz_io_dataIn_1_payload_address_35;
    _zz_io_dataIn_1_payload_address_37 <= _zz_io_dataIn_1_payload_address_36;
    _zz_io_dataIn_1_payload_address_38 <= _zz_io_dataIn_1_payload_address_37;
    _zz_io_dataIn_1_payload_address_39 <= _zz_io_dataIn_1_payload_address_38;
    _zz_io_dataIn_1_payload_address_40 <= _zz_io_dataIn_1_payload_address_39;
    _zz_io_dataIn_1_payload_address_41 <= _zz_io_dataIn_1_payload_address_40;
    _zz_io_dataIn_1_payload_address_42 <= _zz_io_dataIn_1_payload_address_41;
    _zz_io_dataIn_1_payload_address_43 <= _zz_io_dataIn_1_payload_address_42;
    _zz_io_dataIn_1_payload_address_44 <= _zz_io_dataIn_1_payload_address_43;
    _zz_io_dataIn_1_payload_address_45 <= _zz_io_dataIn_1_payload_address_44;
    _zz_io_dataIn_1_payload_address_46 <= _zz_io_dataIn_1_payload_address_45;
    _zz_io_dataIn_1_payload_address_47 <= _zz_io_dataIn_1_payload_address_46;
    _zz_io_dataIn_1_payload_address_48 <= _zz_io_dataIn_1_payload_address_47;
    _zz_io_dataIn_1_payload_address_49 <= _zz_io_dataIn_1_payload_address_48;
    _zz_io_dataIn_1_payload_address_50 <= _zz_io_dataIn_1_payload_address_49;
    _zz_io_dataIn_1_payload_address_51 <= _zz_io_dataIn_1_payload_address_50;
    _zz_io_dataIn_1_payload_address_52 <= _zz_io_dataIn_1_payload_address_51;
    _zz_io_dataIn_1_payload_address_53 <= _zz_io_dataIn_1_payload_address_52;
    _zz_io_dataIn_1_payload_address_54 <= _zz_io_dataIn_1_payload_address_53;
    _zz_io_dataIn_1_payload_address_55 <= _zz_io_dataIn_1_payload_address_54;
    _zz_io_dataIn_1_payload_address_56 <= _zz_io_dataIn_1_payload_address_55;
    _zz_io_dataIn_1_payload_address_57 <= _zz_io_dataIn_1_payload_address_56;
    _zz_io_dataIn_1_payload_address_58 <= _zz_io_dataIn_1_payload_address_57;
    _zz_io_dataIn_1_payload_address_59 <= _zz_io_dataIn_1_payload_address_58;
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      _zz_io_dataIn_1_valid_70 <= 1'b0;
      _zz_io_dataIn_1_valid_71 <= 1'b0;
      _zz_io_dataIn_1_valid_72 <= 1'b0;
      _zz_io_dataIn_1_valid_73 <= 1'b0;
      _zz_io_dataIn_1_valid_74 <= 1'b0;
      _zz_io_dataIn_1_valid_75 <= 1'b0;
      _zz_io_dataIn_1_valid_76 <= 1'b0;
      _zz_io_dataIn_1_valid_77 <= 1'b0;
      _zz_io_dataIn_1_valid_78 <= 1'b0;
      _zz_io_dataIn_1_valid_79 <= 1'b0;
      _zz_io_dataIn_1_valid_80 <= 1'b0;
      _zz_io_dataIn_1_valid_81 <= 1'b0;
      _zz_io_dataIn_1_valid_82 <= 1'b0;
      _zz_io_dataIn_1_valid_83 <= 1'b0;
      _zz_io_dataIn_1_valid_84 <= 1'b0;
      _zz_io_dataIn_1_valid_85 <= 1'b0;
      _zz_io_dataIn_1_valid_86 <= 1'b0;
      _zz_io_dataIn_1_valid_87 <= 1'b0;
      _zz_io_dataIn_1_valid_88 <= 1'b0;
      _zz_io_dataIn_1_valid_89 <= 1'b0;
      _zz_io_dataIn_1_valid_90 <= 1'b0;
      _zz_io_dataIn_1_valid_91 <= 1'b0;
      _zz_io_dataIn_1_valid_92 <= 1'b0;
      _zz_io_dataIn_1_valid_93 <= 1'b0;
      _zz_io_dataIn_1_valid_94 <= 1'b0;
      _zz_io_dataIn_1_valid_95 <= 1'b0;
      _zz_io_dataIn_1_valid_96 <= 1'b0;
      _zz_io_dataIn_1_valid_97 <= 1'b0;
      _zz_io_dataIn_1_valid_98 <= 1'b0;
      _zz_io_dataIn_1_valid_99 <= 1'b0;
      _zz_io_dataIn_1_valid_100 <= 1'b0;
      _zz_io_dataIn_1_valid_101 <= 1'b0;
      _zz_io_dataIn_1_valid_102 <= 1'b0;
      _zz_io_dataIn_1_valid_103 <= 1'b0;
      _zz_io_dataIn_1_valid_104 <= 1'b0;
      _zz_io_dataIn_1_valid_105 <= 1'b0;
      _zz_io_dataIn_1_valid_106 <= 1'b0;
      _zz_io_dataIn_1_valid_107 <= 1'b0;
      _zz_io_dataIn_1_valid_108 <= 1'b0;
      _zz_io_dataIn_1_valid_109 <= 1'b0;
      _zz_io_dataIn_1_valid_110 <= 1'b0;
      _zz_io_dataIn_1_valid_111 <= 1'b0;
      _zz_io_dataIn_1_valid_112 <= 1'b0;
      _zz_io_dataIn_1_valid_113 <= 1'b0;
      _zz_io_dataIn_1_valid_114 <= 1'b0;
      _zz_io_dataIn_1_valid_115 <= 1'b0;
      _zz_io_dataIn_1_valid_116 <= 1'b0;
      _zz_io_dataIn_1_valid_117 <= 1'b0;
      _zz_io_dataIn_1_valid_118 <= 1'b0;
      _zz_io_dataIn_1_valid_119 <= 1'b0;
      _zz_io_dataIn_1_valid_120 <= 1'b0;
      _zz_io_dataIn_1_valid_121 <= 1'b0;
      _zz_io_dataIn_1_valid_122 <= 1'b0;
      _zz_io_dataIn_1_valid_123 <= 1'b0;
      _zz_io_dataIn_1_valid_124 <= 1'b0;
      _zz_io_dataIn_1_valid_125 <= 1'b0;
      _zz_io_dataIn_1_valid_126 <= 1'b0;
      _zz_io_dataIn_1_valid_127 <= 1'b0;
      _zz_io_dataIn_1_valid_128 <= 1'b0;
      _zz_io_dataIn_1_valid_129 <= 1'b0;
    end else begin
      _zz_io_dataIn_1_valid_70 <= (((fsm_stateReg & fsm_enumDef_stage2) != 5'b00000) && (! stage2_calCnt_value[1]));
      _zz_io_dataIn_1_valid_71 <= _zz_io_dataIn_1_valid_70;
      _zz_io_dataIn_1_valid_72 <= _zz_io_dataIn_1_valid_71;
      _zz_io_dataIn_1_valid_73 <= _zz_io_dataIn_1_valid_72;
      _zz_io_dataIn_1_valid_74 <= _zz_io_dataIn_1_valid_73;
      _zz_io_dataIn_1_valid_75 <= _zz_io_dataIn_1_valid_74;
      _zz_io_dataIn_1_valid_76 <= _zz_io_dataIn_1_valid_75;
      _zz_io_dataIn_1_valid_77 <= _zz_io_dataIn_1_valid_76;
      _zz_io_dataIn_1_valid_78 <= _zz_io_dataIn_1_valid_77;
      _zz_io_dataIn_1_valid_79 <= _zz_io_dataIn_1_valid_78;
      _zz_io_dataIn_1_valid_80 <= _zz_io_dataIn_1_valid_79;
      _zz_io_dataIn_1_valid_81 <= _zz_io_dataIn_1_valid_80;
      _zz_io_dataIn_1_valid_82 <= _zz_io_dataIn_1_valid_81;
      _zz_io_dataIn_1_valid_83 <= _zz_io_dataIn_1_valid_82;
      _zz_io_dataIn_1_valid_84 <= _zz_io_dataIn_1_valid_83;
      _zz_io_dataIn_1_valid_85 <= _zz_io_dataIn_1_valid_84;
      _zz_io_dataIn_1_valid_86 <= _zz_io_dataIn_1_valid_85;
      _zz_io_dataIn_1_valid_87 <= _zz_io_dataIn_1_valid_86;
      _zz_io_dataIn_1_valid_88 <= _zz_io_dataIn_1_valid_87;
      _zz_io_dataIn_1_valid_89 <= _zz_io_dataIn_1_valid_88;
      _zz_io_dataIn_1_valid_90 <= _zz_io_dataIn_1_valid_89;
      _zz_io_dataIn_1_valid_91 <= _zz_io_dataIn_1_valid_90;
      _zz_io_dataIn_1_valid_92 <= _zz_io_dataIn_1_valid_91;
      _zz_io_dataIn_1_valid_93 <= _zz_io_dataIn_1_valid_92;
      _zz_io_dataIn_1_valid_94 <= _zz_io_dataIn_1_valid_93;
      _zz_io_dataIn_1_valid_95 <= _zz_io_dataIn_1_valid_94;
      _zz_io_dataIn_1_valid_96 <= _zz_io_dataIn_1_valid_95;
      _zz_io_dataIn_1_valid_97 <= _zz_io_dataIn_1_valid_96;
      _zz_io_dataIn_1_valid_98 <= _zz_io_dataIn_1_valid_97;
      _zz_io_dataIn_1_valid_99 <= _zz_io_dataIn_1_valid_98;
      _zz_io_dataIn_1_valid_100 <= (((fsm_stateReg & fsm_enumDef_stage2) != 5'b00000) && (! stage2_calCnt_value[1]));
      _zz_io_dataIn_1_valid_101 <= _zz_io_dataIn_1_valid_100;
      _zz_io_dataIn_1_valid_102 <= _zz_io_dataIn_1_valid_101;
      _zz_io_dataIn_1_valid_103 <= _zz_io_dataIn_1_valid_102;
      _zz_io_dataIn_1_valid_104 <= _zz_io_dataIn_1_valid_103;
      _zz_io_dataIn_1_valid_105 <= _zz_io_dataIn_1_valid_104;
      _zz_io_dataIn_1_valid_106 <= _zz_io_dataIn_1_valid_105;
      _zz_io_dataIn_1_valid_107 <= _zz_io_dataIn_1_valid_106;
      _zz_io_dataIn_1_valid_108 <= _zz_io_dataIn_1_valid_107;
      _zz_io_dataIn_1_valid_109 <= _zz_io_dataIn_1_valid_108;
      _zz_io_dataIn_1_valid_110 <= _zz_io_dataIn_1_valid_109;
      _zz_io_dataIn_1_valid_111 <= _zz_io_dataIn_1_valid_110;
      _zz_io_dataIn_1_valid_112 <= _zz_io_dataIn_1_valid_111;
      _zz_io_dataIn_1_valid_113 <= _zz_io_dataIn_1_valid_112;
      _zz_io_dataIn_1_valid_114 <= _zz_io_dataIn_1_valid_113;
      _zz_io_dataIn_1_valid_115 <= _zz_io_dataIn_1_valid_114;
      _zz_io_dataIn_1_valid_116 <= _zz_io_dataIn_1_valid_115;
      _zz_io_dataIn_1_valid_117 <= _zz_io_dataIn_1_valid_116;
      _zz_io_dataIn_1_valid_118 <= _zz_io_dataIn_1_valid_117;
      _zz_io_dataIn_1_valid_119 <= _zz_io_dataIn_1_valid_118;
      _zz_io_dataIn_1_valid_120 <= _zz_io_dataIn_1_valid_119;
      _zz_io_dataIn_1_valid_121 <= _zz_io_dataIn_1_valid_120;
      _zz_io_dataIn_1_valid_122 <= _zz_io_dataIn_1_valid_121;
      _zz_io_dataIn_1_valid_123 <= _zz_io_dataIn_1_valid_122;
      _zz_io_dataIn_1_valid_124 <= _zz_io_dataIn_1_valid_123;
      _zz_io_dataIn_1_valid_125 <= _zz_io_dataIn_1_valid_124;
      _zz_io_dataIn_1_valid_126 <= _zz_io_dataIn_1_valid_125;
      _zz_io_dataIn_1_valid_127 <= _zz_io_dataIn_1_valid_126;
      _zz_io_dataIn_1_valid_128 <= _zz_io_dataIn_1_valid_127;
      _zz_io_dataIn_1_valid_129 <= _zz_io_dataIn_1_valid_128;
    end
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      _zz_io_dataIn_1_valid_130 <= 1'b0;
      _zz_io_dataIn_1_valid_131 <= 1'b0;
      _zz_io_dataIn_1_valid_132 <= 1'b0;
      _zz_io_dataIn_1_valid_133 <= 1'b0;
      _zz_io_dataIn_1_valid_134 <= 1'b0;
      _zz_io_dataIn_1_valid_135 <= 1'b0;
      _zz_io_dataIn_1_valid_136 <= 1'b0;
      _zz_io_dataIn_1_valid_137 <= 1'b0;
      _zz_io_dataIn_1_valid_138 <= 1'b0;
      _zz_io_dataIn_1_valid_139 <= 1'b0;
      _zz_io_dataIn_1_valid_140 <= 1'b0;
      _zz_io_dataIn_1_valid_141 <= 1'b0;
      _zz_io_dataIn_1_valid_142 <= 1'b0;
      _zz_io_dataIn_1_valid_143 <= 1'b0;
      _zz_io_dataIn_1_valid_144 <= 1'b0;
      _zz_io_dataIn_1_valid_145 <= 1'b0;
      _zz_io_dataIn_1_valid_146 <= 1'b0;
      _zz_io_dataIn_1_valid_147 <= 1'b0;
      _zz_io_dataIn_1_valid_148 <= 1'b0;
      _zz_io_dataIn_1_valid_149 <= 1'b0;
      _zz_io_dataIn_1_valid_150 <= 1'b0;
      _zz_io_dataIn_1_valid_151 <= 1'b0;
      _zz_io_dataIn_1_valid_152 <= 1'b0;
      _zz_io_dataIn_1_valid_153 <= 1'b0;
      _zz_io_dataIn_1_valid_154 <= 1'b0;
      _zz_io_dataIn_1_valid_155 <= 1'b0;
      _zz_io_dataIn_1_valid_156 <= 1'b0;
      _zz_io_dataIn_1_valid_157 <= 1'b0;
      _zz_io_dataIn_1_valid_158 <= 1'b0;
      _zz_io_dataIn_1_valid_159 <= 1'b0;
      _zz_io_dataIn_1_valid_160 <= 1'b0;
      _zz_io_dataIn_1_valid_161 <= 1'b0;
      _zz_io_dataIn_1_valid_162 <= 1'b0;
      _zz_io_dataIn_1_valid_163 <= 1'b0;
      _zz_io_dataIn_1_valid_164 <= 1'b0;
      _zz_io_dataIn_1_valid_165 <= 1'b0;
      _zz_io_dataIn_1_valid_166 <= 1'b0;
      _zz_io_dataIn_1_valid_167 <= 1'b0;
      _zz_io_dataIn_1_valid_168 <= 1'b0;
      _zz_io_dataIn_1_valid_169 <= 1'b0;
      _zz_io_dataIn_1_valid_170 <= 1'b0;
      _zz_io_dataIn_1_valid_171 <= 1'b0;
      _zz_io_dataIn_1_valid_172 <= 1'b0;
      _zz_io_dataIn_1_valid_173 <= 1'b0;
      _zz_io_dataIn_1_valid_174 <= 1'b0;
      _zz_io_dataIn_1_valid_175 <= 1'b0;
      _zz_io_dataIn_1_valid_176 <= 1'b0;
      _zz_io_dataIn_1_valid_177 <= 1'b0;
      _zz_io_dataIn_1_valid_178 <= 1'b0;
      _zz_io_dataIn_1_valid_179 <= 1'b0;
      _zz_io_dataIn_1_valid_180 <= 1'b0;
      _zz_io_dataIn_1_valid_181 <= 1'b0;
      _zz_io_dataIn_1_valid_182 <= 1'b0;
      _zz_io_dataIn_1_valid_183 <= 1'b0;
      _zz_io_dataIn_1_valid_184 <= 1'b0;
      _zz_io_dataIn_1_valid_185 <= 1'b0;
      _zz_io_dataIn_1_valid_186 <= 1'b0;
      _zz_io_dataIn_1_valid_187 <= 1'b0;
      _zz_io_dataIn_1_valid_188 <= 1'b0;
      _zz_io_dataIn_1_valid_189 <= 1'b0;
    end else begin
      _zz_io_dataIn_1_valid_130 <= ((stage3_doubleWaitCnt_value == 9'h001) || (stage3_addWaitCnt_value == 9'h001));
      _zz_io_dataIn_1_valid_131 <= _zz_io_dataIn_1_valid_130;
      _zz_io_dataIn_1_valid_132 <= _zz_io_dataIn_1_valid_131;
      _zz_io_dataIn_1_valid_133 <= _zz_io_dataIn_1_valid_132;
      _zz_io_dataIn_1_valid_134 <= _zz_io_dataIn_1_valid_133;
      _zz_io_dataIn_1_valid_135 <= _zz_io_dataIn_1_valid_134;
      _zz_io_dataIn_1_valid_136 <= _zz_io_dataIn_1_valid_135;
      _zz_io_dataIn_1_valid_137 <= _zz_io_dataIn_1_valid_136;
      _zz_io_dataIn_1_valid_138 <= _zz_io_dataIn_1_valid_137;
      _zz_io_dataIn_1_valid_139 <= _zz_io_dataIn_1_valid_138;
      _zz_io_dataIn_1_valid_140 <= _zz_io_dataIn_1_valid_139;
      _zz_io_dataIn_1_valid_141 <= _zz_io_dataIn_1_valid_140;
      _zz_io_dataIn_1_valid_142 <= _zz_io_dataIn_1_valid_141;
      _zz_io_dataIn_1_valid_143 <= _zz_io_dataIn_1_valid_142;
      _zz_io_dataIn_1_valid_144 <= _zz_io_dataIn_1_valid_143;
      _zz_io_dataIn_1_valid_145 <= _zz_io_dataIn_1_valid_144;
      _zz_io_dataIn_1_valid_146 <= _zz_io_dataIn_1_valid_145;
      _zz_io_dataIn_1_valid_147 <= _zz_io_dataIn_1_valid_146;
      _zz_io_dataIn_1_valid_148 <= _zz_io_dataIn_1_valid_147;
      _zz_io_dataIn_1_valid_149 <= _zz_io_dataIn_1_valid_148;
      _zz_io_dataIn_1_valid_150 <= _zz_io_dataIn_1_valid_149;
      _zz_io_dataIn_1_valid_151 <= _zz_io_dataIn_1_valid_150;
      _zz_io_dataIn_1_valid_152 <= _zz_io_dataIn_1_valid_151;
      _zz_io_dataIn_1_valid_153 <= _zz_io_dataIn_1_valid_152;
      _zz_io_dataIn_1_valid_154 <= _zz_io_dataIn_1_valid_153;
      _zz_io_dataIn_1_valid_155 <= _zz_io_dataIn_1_valid_154;
      _zz_io_dataIn_1_valid_156 <= _zz_io_dataIn_1_valid_155;
      _zz_io_dataIn_1_valid_157 <= _zz_io_dataIn_1_valid_156;
      _zz_io_dataIn_1_valid_158 <= _zz_io_dataIn_1_valid_157;
      _zz_io_dataIn_1_valid_159 <= _zz_io_dataIn_1_valid_158;
      _zz_io_dataIn_1_valid_160 <= ((stage3_doubleWaitCnt_value == 9'h001) || (stage3_addWaitCnt_value == 9'h001));
      _zz_io_dataIn_1_valid_161 <= _zz_io_dataIn_1_valid_160;
      _zz_io_dataIn_1_valid_162 <= _zz_io_dataIn_1_valid_161;
      _zz_io_dataIn_1_valid_163 <= _zz_io_dataIn_1_valid_162;
      _zz_io_dataIn_1_valid_164 <= _zz_io_dataIn_1_valid_163;
      _zz_io_dataIn_1_valid_165 <= _zz_io_dataIn_1_valid_164;
      _zz_io_dataIn_1_valid_166 <= _zz_io_dataIn_1_valid_165;
      _zz_io_dataIn_1_valid_167 <= _zz_io_dataIn_1_valid_166;
      _zz_io_dataIn_1_valid_168 <= _zz_io_dataIn_1_valid_167;
      _zz_io_dataIn_1_valid_169 <= _zz_io_dataIn_1_valid_168;
      _zz_io_dataIn_1_valid_170 <= _zz_io_dataIn_1_valid_169;
      _zz_io_dataIn_1_valid_171 <= _zz_io_dataIn_1_valid_170;
      _zz_io_dataIn_1_valid_172 <= _zz_io_dataIn_1_valid_171;
      _zz_io_dataIn_1_valid_173 <= _zz_io_dataIn_1_valid_172;
      _zz_io_dataIn_1_valid_174 <= _zz_io_dataIn_1_valid_173;
      _zz_io_dataIn_1_valid_175 <= _zz_io_dataIn_1_valid_174;
      _zz_io_dataIn_1_valid_176 <= _zz_io_dataIn_1_valid_175;
      _zz_io_dataIn_1_valid_177 <= _zz_io_dataIn_1_valid_176;
      _zz_io_dataIn_1_valid_178 <= _zz_io_dataIn_1_valid_177;
      _zz_io_dataIn_1_valid_179 <= _zz_io_dataIn_1_valid_178;
      _zz_io_dataIn_1_valid_180 <= _zz_io_dataIn_1_valid_179;
      _zz_io_dataIn_1_valid_181 <= _zz_io_dataIn_1_valid_180;
      _zz_io_dataIn_1_valid_182 <= _zz_io_dataIn_1_valid_181;
      _zz_io_dataIn_1_valid_183 <= _zz_io_dataIn_1_valid_182;
      _zz_io_dataIn_1_valid_184 <= _zz_io_dataIn_1_valid_183;
      _zz_io_dataIn_1_valid_185 <= _zz_io_dataIn_1_valid_184;
      _zz_io_dataIn_1_valid_186 <= _zz_io_dataIn_1_valid_185;
      _zz_io_dataIn_1_valid_187 <= _zz_io_dataIn_1_valid_186;
      _zz_io_dataIn_1_valid_188 <= _zz_io_dataIn_1_valid_187;
      _zz_io_dataIn_1_valid_189 <= _zz_io_dataIn_1_valid_188;
    end
  end

  always @(posedge clk) begin
    pippenger_1_dataRam_0_io_rData_1_regNext_X_1 <= dataRam_0_io_rData_1_X;
    pippenger_1_dataRam_0_io_rData_1_regNext_Y_1 <= dataRam_0_io_rData_1_Y;
    pippenger_1_dataRam_0_io_rData_1_regNext_Z_1 <= dataRam_0_io_rData_1_Z;
    pippenger_1_dataRam_0_io_rData_1_regNext_T_1 <= dataRam_0_io_rData_1_T;
    _zz_io_dataIn_1_payload_address_60 <= (stage3_GCnt_value - _zz__zz_io_dataIn_1_payload_address_60);
    _zz_io_dataIn_1_payload_address_61 <= _zz_io_dataIn_1_payload_address_60;
    _zz_io_dataIn_1_payload_address_62 <= _zz_io_dataIn_1_payload_address_61;
    _zz_io_dataIn_1_payload_address_63 <= _zz_io_dataIn_1_payload_address_62;
    _zz_io_dataIn_1_payload_address_64 <= _zz_io_dataIn_1_payload_address_63;
    _zz_io_dataIn_1_payload_address_65 <= _zz_io_dataIn_1_payload_address_64;
    _zz_io_dataIn_1_payload_address_66 <= _zz_io_dataIn_1_payload_address_65;
    _zz_io_dataIn_1_payload_address_67 <= _zz_io_dataIn_1_payload_address_66;
    _zz_io_dataIn_1_payload_address_68 <= _zz_io_dataIn_1_payload_address_67;
    _zz_io_dataIn_1_payload_address_69 <= _zz_io_dataIn_1_payload_address_68;
    _zz_io_dataIn_1_payload_address_70 <= _zz_io_dataIn_1_payload_address_69;
    _zz_io_dataIn_1_payload_address_71 <= _zz_io_dataIn_1_payload_address_70;
    _zz_io_dataIn_1_payload_address_72 <= _zz_io_dataIn_1_payload_address_71;
    _zz_io_dataIn_1_payload_address_73 <= _zz_io_dataIn_1_payload_address_72;
    _zz_io_dataIn_1_payload_address_74 <= _zz_io_dataIn_1_payload_address_73;
    _zz_io_dataIn_1_payload_address_75 <= _zz_io_dataIn_1_payload_address_74;
    _zz_io_dataIn_1_payload_address_76 <= _zz_io_dataIn_1_payload_address_75;
    _zz_io_dataIn_1_payload_address_77 <= _zz_io_dataIn_1_payload_address_76;
    _zz_io_dataIn_1_payload_address_78 <= _zz_io_dataIn_1_payload_address_77;
    _zz_io_dataIn_1_payload_address_79 <= _zz_io_dataIn_1_payload_address_78;
    _zz_io_dataIn_1_payload_address_80 <= _zz_io_dataIn_1_payload_address_79;
    _zz_io_dataIn_1_payload_address_81 <= _zz_io_dataIn_1_payload_address_80;
    _zz_io_dataIn_1_payload_address_82 <= _zz_io_dataIn_1_payload_address_81;
    _zz_io_dataIn_1_payload_address_83 <= _zz_io_dataIn_1_payload_address_82;
    _zz_io_dataIn_1_payload_address_84 <= _zz_io_dataIn_1_payload_address_83;
    _zz_io_dataIn_1_payload_address_85 <= _zz_io_dataIn_1_payload_address_84;
    _zz_io_dataIn_1_payload_address_86 <= _zz_io_dataIn_1_payload_address_85;
    _zz_io_dataIn_1_payload_address_87 <= _zz_io_dataIn_1_payload_address_86;
    _zz_io_dataIn_1_payload_address_88 <= _zz_io_dataIn_1_payload_address_87;
    _zz_io_dataIn_1_payload_address_89 <= _zz_io_dataIn_1_payload_address_88;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_X_1 <= dataRam_1_1_io_rData_1_X;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_1 <= dataRam_1_1_io_rData_1_Y;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_1 <= dataRam_1_1_io_rData_1_Z;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_T_1 <= dataRam_1_1_io_rData_1_T;
    _zz_io_dataIn_1_payload_address_90 <= (stage3_GCnt_value - _zz__zz_io_dataIn_1_payload_address_90);
    _zz_io_dataIn_1_payload_address_91 <= _zz_io_dataIn_1_payload_address_90;
    _zz_io_dataIn_1_payload_address_92 <= _zz_io_dataIn_1_payload_address_91;
    _zz_io_dataIn_1_payload_address_93 <= _zz_io_dataIn_1_payload_address_92;
    _zz_io_dataIn_1_payload_address_94 <= _zz_io_dataIn_1_payload_address_93;
    _zz_io_dataIn_1_payload_address_95 <= _zz_io_dataIn_1_payload_address_94;
    _zz_io_dataIn_1_payload_address_96 <= _zz_io_dataIn_1_payload_address_95;
    _zz_io_dataIn_1_payload_address_97 <= _zz_io_dataIn_1_payload_address_96;
    _zz_io_dataIn_1_payload_address_98 <= _zz_io_dataIn_1_payload_address_97;
    _zz_io_dataIn_1_payload_address_99 <= _zz_io_dataIn_1_payload_address_98;
    _zz_io_dataIn_1_payload_address_100 <= _zz_io_dataIn_1_payload_address_99;
    _zz_io_dataIn_1_payload_address_101 <= _zz_io_dataIn_1_payload_address_100;
    _zz_io_dataIn_1_payload_address_102 <= _zz_io_dataIn_1_payload_address_101;
    _zz_io_dataIn_1_payload_address_103 <= _zz_io_dataIn_1_payload_address_102;
    _zz_io_dataIn_1_payload_address_104 <= _zz_io_dataIn_1_payload_address_103;
    _zz_io_dataIn_1_payload_address_105 <= _zz_io_dataIn_1_payload_address_104;
    _zz_io_dataIn_1_payload_address_106 <= _zz_io_dataIn_1_payload_address_105;
    _zz_io_dataIn_1_payload_address_107 <= _zz_io_dataIn_1_payload_address_106;
    _zz_io_dataIn_1_payload_address_108 <= _zz_io_dataIn_1_payload_address_107;
    _zz_io_dataIn_1_payload_address_109 <= _zz_io_dataIn_1_payload_address_108;
    _zz_io_dataIn_1_payload_address_110 <= _zz_io_dataIn_1_payload_address_109;
    _zz_io_dataIn_1_payload_address_111 <= _zz_io_dataIn_1_payload_address_110;
    _zz_io_dataIn_1_payload_address_112 <= _zz_io_dataIn_1_payload_address_111;
    _zz_io_dataIn_1_payload_address_113 <= _zz_io_dataIn_1_payload_address_112;
    _zz_io_dataIn_1_payload_address_114 <= _zz_io_dataIn_1_payload_address_113;
    _zz_io_dataIn_1_payload_address_115 <= _zz_io_dataIn_1_payload_address_114;
    _zz_io_dataIn_1_payload_address_116 <= _zz_io_dataIn_1_payload_address_115;
    _zz_io_dataIn_1_payload_address_117 <= _zz_io_dataIn_1_payload_address_116;
    _zz_io_dataIn_1_payload_address_118 <= _zz_io_dataIn_1_payload_address_117;
    _zz_io_dataIn_1_payload_address_119 <= _zz_io_dataIn_1_payload_address_118;
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      _zz_io_dataIn_1_valid_190 <= 1'b0;
      _zz_io_dataIn_1_valid_191 <= 1'b0;
      _zz_io_dataIn_1_valid_192 <= 1'b0;
      _zz_io_dataIn_1_valid_193 <= 1'b0;
      _zz_io_dataIn_1_valid_194 <= 1'b0;
      _zz_io_dataIn_1_valid_195 <= 1'b0;
      _zz_io_dataIn_1_valid_196 <= 1'b0;
      _zz_io_dataIn_1_valid_197 <= 1'b0;
      _zz_io_dataIn_1_valid_198 <= 1'b0;
      _zz_io_dataIn_1_valid_199 <= 1'b0;
      _zz_io_dataIn_1_valid_200 <= 1'b0;
      _zz_io_dataIn_1_valid_201 <= 1'b0;
      _zz_io_dataIn_1_valid_202 <= 1'b0;
      _zz_io_dataIn_1_valid_203 <= 1'b0;
      _zz_io_dataIn_1_valid_204 <= 1'b0;
      _zz_io_dataIn_1_valid_205 <= 1'b0;
      _zz_io_dataIn_1_valid_206 <= 1'b0;
      _zz_io_dataIn_1_valid_207 <= 1'b0;
      _zz_io_dataIn_1_valid_208 <= 1'b0;
      _zz_io_dataIn_1_valid_209 <= 1'b0;
      _zz_io_dataIn_1_valid_210 <= 1'b0;
      _zz_io_dataIn_1_valid_211 <= 1'b0;
      _zz_io_dataIn_1_valid_212 <= 1'b0;
      _zz_io_dataIn_1_valid_213 <= 1'b0;
      _zz_io_dataIn_1_valid_214 <= 1'b0;
      _zz_io_dataIn_1_valid_215 <= 1'b0;
      _zz_io_dataIn_1_valid_216 <= 1'b0;
      _zz_io_dataIn_1_valid_217 <= 1'b0;
      _zz_io_dataIn_1_valid_218 <= 1'b0;
      _zz_io_dataIn_1_valid_219 <= 1'b0;
      _zz_io_dataIn_1_valid_220 <= 1'b0;
      _zz_io_dataIn_1_valid_221 <= 1'b0;
      _zz_io_dataIn_1_valid_222 <= 1'b0;
      _zz_io_dataIn_1_valid_223 <= 1'b0;
      _zz_io_dataIn_1_valid_224 <= 1'b0;
      _zz_io_dataIn_1_valid_225 <= 1'b0;
      _zz_io_dataIn_1_valid_226 <= 1'b0;
      _zz_io_dataIn_1_valid_227 <= 1'b0;
      _zz_io_dataIn_1_valid_228 <= 1'b0;
      _zz_io_dataIn_1_valid_229 <= 1'b0;
      _zz_io_dataIn_1_valid_230 <= 1'b0;
      _zz_io_dataIn_1_valid_231 <= 1'b0;
      _zz_io_dataIn_1_valid_232 <= 1'b0;
      _zz_io_dataIn_1_valid_233 <= 1'b0;
      _zz_io_dataIn_1_valid_234 <= 1'b0;
      _zz_io_dataIn_1_valid_235 <= 1'b0;
      _zz_io_dataIn_1_valid_236 <= 1'b0;
      _zz_io_dataIn_1_valid_237 <= 1'b0;
      _zz_io_dataIn_1_valid_238 <= 1'b0;
      _zz_io_dataIn_1_valid_239 <= 1'b0;
      _zz_io_dataIn_1_valid_240 <= 1'b0;
      _zz_io_dataIn_1_valid_241 <= 1'b0;
      _zz_io_dataIn_1_valid_242 <= 1'b0;
      _zz_io_dataIn_1_valid_243 <= 1'b0;
      _zz_io_dataIn_1_valid_244 <= 1'b0;
      _zz_io_dataIn_1_valid_245 <= 1'b0;
      _zz_io_dataIn_1_valid_246 <= 1'b0;
      _zz_io_dataIn_1_valid_247 <= 1'b0;
      _zz_io_dataIn_1_valid_248 <= 1'b0;
      _zz_io_dataIn_1_valid_249 <= 1'b0;
    end else begin
      _zz_io_dataIn_1_valid_190 <= ((stage3Final_addWaitCnt_value == 9'h001) && stage3Final_pAddShr[0]);
      _zz_io_dataIn_1_valid_191 <= _zz_io_dataIn_1_valid_190;
      _zz_io_dataIn_1_valid_192 <= _zz_io_dataIn_1_valid_191;
      _zz_io_dataIn_1_valid_193 <= _zz_io_dataIn_1_valid_192;
      _zz_io_dataIn_1_valid_194 <= _zz_io_dataIn_1_valid_193;
      _zz_io_dataIn_1_valid_195 <= _zz_io_dataIn_1_valid_194;
      _zz_io_dataIn_1_valid_196 <= _zz_io_dataIn_1_valid_195;
      _zz_io_dataIn_1_valid_197 <= _zz_io_dataIn_1_valid_196;
      _zz_io_dataIn_1_valid_198 <= _zz_io_dataIn_1_valid_197;
      _zz_io_dataIn_1_valid_199 <= _zz_io_dataIn_1_valid_198;
      _zz_io_dataIn_1_valid_200 <= _zz_io_dataIn_1_valid_199;
      _zz_io_dataIn_1_valid_201 <= _zz_io_dataIn_1_valid_200;
      _zz_io_dataIn_1_valid_202 <= _zz_io_dataIn_1_valid_201;
      _zz_io_dataIn_1_valid_203 <= _zz_io_dataIn_1_valid_202;
      _zz_io_dataIn_1_valid_204 <= _zz_io_dataIn_1_valid_203;
      _zz_io_dataIn_1_valid_205 <= _zz_io_dataIn_1_valid_204;
      _zz_io_dataIn_1_valid_206 <= _zz_io_dataIn_1_valid_205;
      _zz_io_dataIn_1_valid_207 <= _zz_io_dataIn_1_valid_206;
      _zz_io_dataIn_1_valid_208 <= _zz_io_dataIn_1_valid_207;
      _zz_io_dataIn_1_valid_209 <= _zz_io_dataIn_1_valid_208;
      _zz_io_dataIn_1_valid_210 <= _zz_io_dataIn_1_valid_209;
      _zz_io_dataIn_1_valid_211 <= _zz_io_dataIn_1_valid_210;
      _zz_io_dataIn_1_valid_212 <= _zz_io_dataIn_1_valid_211;
      _zz_io_dataIn_1_valid_213 <= _zz_io_dataIn_1_valid_212;
      _zz_io_dataIn_1_valid_214 <= _zz_io_dataIn_1_valid_213;
      _zz_io_dataIn_1_valid_215 <= _zz_io_dataIn_1_valid_214;
      _zz_io_dataIn_1_valid_216 <= _zz_io_dataIn_1_valid_215;
      _zz_io_dataIn_1_valid_217 <= _zz_io_dataIn_1_valid_216;
      _zz_io_dataIn_1_valid_218 <= _zz_io_dataIn_1_valid_217;
      _zz_io_dataIn_1_valid_219 <= _zz_io_dataIn_1_valid_218;
      _zz_io_dataIn_1_valid_220 <= ((stage3Final_doubleWaitCnt_value == 9'h001) && stage3Final_pAddShr[0]);
      _zz_io_dataIn_1_valid_221 <= _zz_io_dataIn_1_valid_220;
      _zz_io_dataIn_1_valid_222 <= _zz_io_dataIn_1_valid_221;
      _zz_io_dataIn_1_valid_223 <= _zz_io_dataIn_1_valid_222;
      _zz_io_dataIn_1_valid_224 <= _zz_io_dataIn_1_valid_223;
      _zz_io_dataIn_1_valid_225 <= _zz_io_dataIn_1_valid_224;
      _zz_io_dataIn_1_valid_226 <= _zz_io_dataIn_1_valid_225;
      _zz_io_dataIn_1_valid_227 <= _zz_io_dataIn_1_valid_226;
      _zz_io_dataIn_1_valid_228 <= _zz_io_dataIn_1_valid_227;
      _zz_io_dataIn_1_valid_229 <= _zz_io_dataIn_1_valid_228;
      _zz_io_dataIn_1_valid_230 <= _zz_io_dataIn_1_valid_229;
      _zz_io_dataIn_1_valid_231 <= _zz_io_dataIn_1_valid_230;
      _zz_io_dataIn_1_valid_232 <= _zz_io_dataIn_1_valid_231;
      _zz_io_dataIn_1_valid_233 <= _zz_io_dataIn_1_valid_232;
      _zz_io_dataIn_1_valid_234 <= _zz_io_dataIn_1_valid_233;
      _zz_io_dataIn_1_valid_235 <= _zz_io_dataIn_1_valid_234;
      _zz_io_dataIn_1_valid_236 <= _zz_io_dataIn_1_valid_235;
      _zz_io_dataIn_1_valid_237 <= _zz_io_dataIn_1_valid_236;
      _zz_io_dataIn_1_valid_238 <= _zz_io_dataIn_1_valid_237;
      _zz_io_dataIn_1_valid_239 <= _zz_io_dataIn_1_valid_238;
      _zz_io_dataIn_1_valid_240 <= _zz_io_dataIn_1_valid_239;
      _zz_io_dataIn_1_valid_241 <= _zz_io_dataIn_1_valid_240;
      _zz_io_dataIn_1_valid_242 <= _zz_io_dataIn_1_valid_241;
      _zz_io_dataIn_1_valid_243 <= _zz_io_dataIn_1_valid_242;
      _zz_io_dataIn_1_valid_244 <= _zz_io_dataIn_1_valid_243;
      _zz_io_dataIn_1_valid_245 <= _zz_io_dataIn_1_valid_244;
      _zz_io_dataIn_1_valid_246 <= _zz_io_dataIn_1_valid_245;
      _zz_io_dataIn_1_valid_247 <= _zz_io_dataIn_1_valid_246;
      _zz_io_dataIn_1_valid_248 <= _zz_io_dataIn_1_valid_247;
      _zz_io_dataIn_1_valid_249 <= _zz_io_dataIn_1_valid_248;
    end
  end

  always @(posedge clk) begin
    pippenger_1_dataRam_1_1_io_rData_1_regNext_X_2 <= dataRam_1_1_io_rData_1_X;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_2 <= dataRam_1_1_io_rData_1_Y;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_2 <= dataRam_1_1_io_rData_1_Z;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_T_2 <= dataRam_1_1_io_rData_1_T;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_X_3 <= dataRam_1_1_io_rData_1_X;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_Y_3 <= dataRam_1_1_io_rData_1_Y;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_Z_3 <= dataRam_1_1_io_rData_1_Z;
    pippenger_1_dataRam_1_1_io_rData_1_regNext_T_3 <= dataRam_1_1_io_rData_1_T;
  end


endmodule

module PNeg (
  input      [376:0]  io_a_X,
  input      [376:0]  io_a_Y,
  input      [376:0]  io_a_Z,
  input      [376:0]  io_a_T,
  output     [376:0]  io_n_X,
  output     [376:0]  io_n_Y,
  output     [376:0]  io_n_Z,
  output     [376:0]  io_n_T,
  input               clk,
  input               resetn
);

  wire       [377:0]  sub_io_s;
  reg        [376:0]  io_a_X_delay_1;
  reg        [376:0]  io_a_X_delay_2;
  reg        [376:0]  io_a_X_delay_3;
  reg        [376:0]  io_a_X_delay_4;
  reg        [376:0]  io_a_X_delay_5;
  reg        [376:0]  io_a_X_delay_6;
  reg        [376:0]  io_a_T_delay_1;
  reg        [376:0]  io_a_T_delay_2;
  reg        [376:0]  io_a_T_delay_3;
  reg        [376:0]  io_a_T_delay_4;
  reg        [376:0]  io_a_T_delay_5;
  reg        [376:0]  io_a_T_delay_6;

  BADD sub (
    .io_a   (377'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001), //i
    .io_b   (io_a_Y[376:0]                                                                                       ), //i
    .io_c   (1'b1                                                                                                ), //i
    .io_s   (sub_io_s[377:0]                                                                                     ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  assign io_n_X = io_a_X_delay_6;
  assign io_n_Y = sub_io_s[376:0];
  assign io_n_Z = 377'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000000;
  assign io_n_T = io_a_T_delay_6;
  always @(posedge clk) begin
    io_a_X_delay_1 <= io_a_X;
    io_a_X_delay_2 <= io_a_X_delay_1;
    io_a_X_delay_3 <= io_a_X_delay_2;
    io_a_X_delay_4 <= io_a_X_delay_3;
    io_a_X_delay_5 <= io_a_X_delay_4;
    io_a_X_delay_6 <= io_a_X_delay_5;
    io_a_T_delay_1 <= io_a_T;
    io_a_T_delay_2 <= io_a_T_delay_1;
    io_a_T_delay_3 <= io_a_T_delay_2;
    io_a_T_delay_4 <= io_a_T_delay_3;
    io_a_T_delay_5 <= io_a_T_delay_4;
    io_a_T_delay_6 <= io_a_T_delay_5;
  end


endmodule

module PAdd_1 (
  input      [376:0]  io_a_X,
  input      [376:0]  io_a_Y,
  input      [376:0]  io_a_Z,
  input      [376:0]  io_a_T,
  input      [376:0]  io_b_X,
  input      [376:0]  io_b_Y,
  input      [376:0]  io_b_Z,
  input      [376:0]  io_b_T,
  output     [376:0]  io_s_X,
  output     [376:0]  io_s_Y,
  output     [376:0]  io_s_Z,
  output     [376:0]  io_s_T,
  input               clk,
  input               resetn
);

  wire       [377:0]  reduction_io_a;
  wire       [376:0]  mul_0_io_p;
  wire       [376:0]  mul_1_io_p;
  wire       [376:0]  mul_2_io_p;
  wire       [376:0]  mul_3_io_p;
  wire       [376:0]  mul_4_io_p;
  wire       [376:0]  mul_5_io_p;
  wire       [376:0]  mul_6_io_p;
  wire       [376:0]  mul_7_io_p;
  wire       [376:0]  cMul_io_p;
  wire       [376:0]  add_0_io_s;
  wire       [376:0]  add_1_1_io_s;
  wire       [376:0]  add_2_1_io_s;
  wire       [376:0]  add_3_1_io_s;
  wire       [376:0]  sub_0_io_s;
  wire       [376:0]  sub_1_io_s;
  wire       [376:0]  sub_2_io_s;
  wire       [376:0]  sub_3_io_s;
  wire       [376:0]  reduction_io_r;
  reg        [376:0]  io_a_T_delay_1;
  reg        [376:0]  io_a_T_delay_2;
  reg        [376:0]  io_a_T_delay_3;
  reg        [376:0]  io_a_T_delay_4;
  reg        [376:0]  io_a_T_delay_5;
  reg        [376:0]  io_a_T_delay_6;
  reg        [376:0]  io_a_T_delay_7;
  reg        [376:0]  io_a_T_delay_8;
  reg        [376:0]  io_a_T_delay_9;
  reg        [376:0]  io_a_T_delay_10;
  reg        [376:0]  io_a_T_delay_11;
  reg        [376:0]  io_a_T_delay_12;
  reg        [376:0]  io_a_T_delay_13;
  reg        [376:0]  io_a_T_delay_14;
  reg        [376:0]  io_a_T_delay_15;
  reg        [376:0]  io_a_T_delay_16;
  reg        [376:0]  io_a_T_delay_17;
  reg        [376:0]  io_a_T_delay_18;
  reg        [376:0]  io_a_T_delay_19;
  reg        [376:0]  io_a_T_delay_20;
  reg        [376:0]  io_a_T_delay_21;
  reg        [376:0]  io_a_T_delay_22;
  reg        [376:0]  io_a_T_delay_23;
  reg        [376:0]  io_a_T_delay_24;
  reg        [376:0]  io_a_T_delay_25;
  reg        [376:0]  io_a_T_delay_26;
  reg        [376:0]  io_a_T_delay_27;
  reg        [376:0]  io_a_T_delay_28;
  reg        [376:0]  io_a_T_delay_29;
  reg        [376:0]  io_a_T_delay_30;
  reg        [376:0]  io_a_T_delay_31;
  reg        [376:0]  io_a_T_delay_32;
  reg        [376:0]  io_a_T_delay_33;
  reg        [376:0]  io_a_T_delay_34;
  reg        [376:0]  io_a_T_delay_35;
  reg        [376:0]  io_a_T_delay_36;
  reg        [376:0]  io_a_T_delay_37;
  reg        [376:0]  io_a_T_delay_38;
  reg        [376:0]  io_a_T_delay_39;
  reg        [376:0]  io_a_T_delay_40;
  reg        [376:0]  io_a_T_delay_41;
  reg        [376:0]  io_a_T_delay_42;
  reg        [376:0]  io_a_T_delay_43;
  reg        [376:0]  io_a_T_delay_44;
  reg        [376:0]  io_a_T_delay_45;
  reg        [376:0]  io_a_T_delay_46;
  reg        [376:0]  io_a_T_delay_47;
  reg        [376:0]  io_a_T_delay_48;
  reg        [376:0]  io_a_T_delay_49;
  reg        [376:0]  io_a_T_delay_50;
  reg        [376:0]  io_a_T_delay_51;
  reg        [376:0]  io_a_T_delay_52;
  reg        [376:0]  io_a_T_delay_53;
  reg        [376:0]  io_a_T_delay_54;
  reg        [376:0]  io_a_T_delay_55;
  reg        [376:0]  io_a_T_delay_56;
  reg        [376:0]  io_a_T_delay_57;
  reg        [376:0]  io_a_T_delay_58;
  reg        [376:0]  io_a_T_delay_59;
  reg        [376:0]  io_a_T_delay_60;
  reg        [376:0]  io_a_T_delay_61;
  reg        [376:0]  io_a_T_delay_62;
  reg        [376:0]  io_a_T_delay_63;
  reg        [376:0]  io_a_T_delay_64;
  reg        [376:0]  io_a_T_delay_65;
  reg        [376:0]  io_a_T_delay_66;
  reg        [376:0]  io_a_T_delay_67;
  reg        [376:0]  io_a_T_delay_68;
  reg        [376:0]  io_a_T_delay_69;
  reg        [376:0]  io_a_T_delay_70;
  reg        [376:0]  io_a_T_delay_71;
  reg        [376:0]  io_a_T_delay_72;
  reg        [376:0]  io_a_T_delay_73;
  reg        [376:0]  io_a_T_delay_74;
  reg        [376:0]  io_a_T_delay_75;
  reg        [376:0]  io_a_T_delay_76;
  reg        [376:0]  io_a_T_delay_77;
  reg        [376:0]  io_a_T_delay_78;
  reg        [376:0]  io_a_T_delay_79;
  reg        [376:0]  io_a_T_delay_80;
  reg        [376:0]  io_a_T_delay_81;
  reg        [376:0]  io_a_T_delay_82;
  reg        [376:0]  io_a_T_delay_83;
  reg        [376:0]  io_a_T_delay_84;
  reg        [376:0]  adder_1_reduction_io_r_delay_1;
  reg        [376:0]  adder_1_reduction_io_r_delay_2;
  reg        [376:0]  adder_1_reduction_io_r_delay_3;
  reg        [376:0]  adder_1_reduction_io_r_delay_4;
  reg        [376:0]  adder_1_reduction_io_r_delay_5;
  reg        [376:0]  adder_1_reduction_io_r_delay_6;
  reg        [376:0]  adder_1_reduction_io_r_delay_7;
  reg        [376:0]  adder_1_reduction_io_r_delay_8;
  reg        [376:0]  adder_1_reduction_io_r_delay_9;
  reg        [376:0]  adder_1_reduction_io_r_delay_10;
  reg        [376:0]  adder_1_reduction_io_r_delay_11;
  reg        [376:0]  adder_1_reduction_io_r_delay_12;
  reg        [376:0]  adder_1_reduction_io_r_delay_13;
  reg        [376:0]  adder_1_reduction_io_r_delay_14;
  reg        [376:0]  adder_1_reduction_io_r_delay_15;
  reg        [376:0]  adder_1_reduction_io_r_delay_16;
  reg        [376:0]  adder_1_reduction_io_r_delay_17;
  reg        [376:0]  adder_1_reduction_io_r_delay_18;
  reg        [376:0]  adder_1_reduction_io_r_delay_19;
  reg        [376:0]  adder_1_reduction_io_r_delay_20;
  reg        [376:0]  adder_1_reduction_io_r_delay_21;
  reg        [376:0]  adder_1_reduction_io_r_delay_22;
  reg        [376:0]  adder_1_reduction_io_r_delay_23;
  reg        [376:0]  adder_1_reduction_io_r_delay_24;
  reg        [376:0]  adder_1_reduction_io_r_delay_25;
  reg        [376:0]  adder_1_reduction_io_r_delay_26;
  reg        [376:0]  adder_1_reduction_io_r_delay_27;
  reg        [376:0]  adder_1_reduction_io_r_delay_28;
  reg        [376:0]  adder_1_reduction_io_r_delay_29;
  reg        [376:0]  adder_1_reduction_io_r_delay_30;
  reg        [376:0]  adder_1_reduction_io_r_delay_31;
  reg        [376:0]  adder_1_reduction_io_r_delay_32;
  reg        [376:0]  adder_1_reduction_io_r_delay_33;
  reg        [376:0]  adder_1_reduction_io_r_delay_34;
  reg        [376:0]  adder_1_reduction_io_r_delay_35;
  reg        [376:0]  adder_1_reduction_io_r_delay_36;
  reg        [376:0]  adder_1_reduction_io_r_delay_37;
  reg        [376:0]  adder_1_reduction_io_r_delay_38;
  reg        [376:0]  adder_1_reduction_io_r_delay_39;
  reg        [376:0]  adder_1_reduction_io_r_delay_40;
  reg        [376:0]  adder_1_reduction_io_r_delay_41;
  reg        [376:0]  adder_1_reduction_io_r_delay_42;
  reg        [376:0]  adder_1_reduction_io_r_delay_43;
  reg        [376:0]  adder_1_reduction_io_r_delay_44;
  reg        [376:0]  adder_1_reduction_io_r_delay_45;
  reg        [376:0]  adder_1_reduction_io_r_delay_46;
  reg        [376:0]  adder_1_reduction_io_r_delay_47;
  reg        [376:0]  adder_1_reduction_io_r_delay_48;
  reg        [376:0]  adder_1_reduction_io_r_delay_49;
  reg        [376:0]  adder_1_reduction_io_r_delay_50;
  reg        [376:0]  adder_1_reduction_io_r_delay_51;
  reg        [376:0]  adder_1_reduction_io_r_delay_52;
  reg        [376:0]  adder_1_reduction_io_r_delay_53;
  reg        [376:0]  adder_1_reduction_io_r_delay_54;
  reg        [376:0]  adder_1_reduction_io_r_delay_55;
  reg        [376:0]  adder_1_reduction_io_r_delay_56;
  reg        [376:0]  adder_1_reduction_io_r_delay_57;
  reg        [376:0]  adder_1_reduction_io_r_delay_58;
  reg        [376:0]  adder_1_reduction_io_r_delay_59;
  reg        [376:0]  adder_1_reduction_io_r_delay_60;
  reg        [376:0]  adder_1_reduction_io_r_delay_61;
  reg        [376:0]  adder_1_reduction_io_r_delay_62;
  reg        [376:0]  adder_1_reduction_io_r_delay_63;
  reg        [376:0]  adder_1_reduction_io_r_delay_64;
  reg        [376:0]  adder_1_reduction_io_r_delay_65;
  reg        [376:0]  adder_1_reduction_io_r_delay_66;
  reg        [376:0]  adder_1_reduction_io_r_delay_67;
  reg        [376:0]  adder_1_reduction_io_r_delay_68;
  reg        [376:0]  adder_1_reduction_io_r_delay_69;
  reg        [376:0]  adder_1_reduction_io_r_delay_70;
  reg        [376:0]  adder_1_reduction_io_r_delay_71;
  reg        [376:0]  adder_1_reduction_io_r_delay_72;
  reg        [376:0]  adder_1_reduction_io_r_delay_73;
  reg        [376:0]  adder_1_reduction_io_r_delay_74;
  reg        [376:0]  adder_1_reduction_io_r_delay_75;
  reg        [376:0]  adder_1_reduction_io_r_delay_76;
  reg        [376:0]  R8;
  reg        [376:0]  adder_1_sub_2_io_s_delay_1;
  reg        [376:0]  adder_1_sub_2_io_s_delay_2;
  reg        [376:0]  adder_1_sub_2_io_s_delay_3;
  reg        [376:0]  adder_1_sub_2_io_s_delay_4;
  reg        [376:0]  adder_1_sub_2_io_s_delay_5;
  reg        [376:0]  adder_1_sub_2_io_s_delay_6;
  reg        [376:0]  adder_1_sub_2_io_s_delay_7;
  reg        [376:0]  adder_1_sub_2_io_s_delay_8;
  reg        [376:0]  adder_1_sub_2_io_s_delay_9;
  reg        [376:0]  adder_1_sub_2_io_s_delay_10;
  reg        [376:0]  adder_1_sub_2_io_s_delay_11;
  reg        [376:0]  adder_1_sub_2_io_s_delay_12;
  reg        [376:0]  adder_1_sub_2_io_s_delay_13;
  reg        [376:0]  adder_1_sub_2_io_s_delay_14;
  reg        [376:0]  adder_1_sub_2_io_s_delay_15;
  reg        [376:0]  adder_1_sub_2_io_s_delay_16;
  reg        [376:0]  adder_1_sub_2_io_s_delay_17;
  reg        [376:0]  adder_1_sub_2_io_s_delay_18;
  reg        [376:0]  adder_1_sub_2_io_s_delay_19;
  reg        [376:0]  adder_1_sub_2_io_s_delay_20;
  reg        [376:0]  adder_1_sub_2_io_s_delay_21;
  reg        [376:0]  adder_1_sub_2_io_s_delay_22;
  reg        [376:0]  adder_1_sub_2_io_s_delay_23;
  reg        [376:0]  adder_1_sub_2_io_s_delay_24;
  reg        [376:0]  adder_1_sub_2_io_s_delay_25;
  reg        [376:0]  adder_1_sub_2_io_s_delay_26;
  reg        [376:0]  adder_1_sub_2_io_s_delay_27;
  reg        [376:0]  adder_1_sub_2_io_s_delay_28;
  reg        [376:0]  adder_1_sub_2_io_s_delay_29;
  reg        [376:0]  adder_1_sub_2_io_s_delay_30;
  reg        [376:0]  adder_1_sub_2_io_s_delay_31;
  reg        [376:0]  adder_1_sub_2_io_s_delay_32;
  reg        [376:0]  adder_1_sub_2_io_s_delay_33;
  reg        [376:0]  adder_1_sub_2_io_s_delay_34;
  reg        [376:0]  adder_1_sub_2_io_s_delay_35;
  reg        [376:0]  adder_1_sub_2_io_s_delay_36;
  reg        [376:0]  adder_1_sub_2_io_s_delay_37;
  reg        [376:0]  adder_1_sub_2_io_s_delay_38;
  reg        [376:0]  adder_1_sub_2_io_s_delay_39;
  reg        [376:0]  adder_1_sub_2_io_s_delay_40;
  reg        [376:0]  adder_1_sub_2_io_s_delay_41;
  reg        [376:0]  adder_1_sub_2_io_s_delay_42;
  reg        [376:0]  adder_1_sub_2_io_s_delay_43;
  reg        [376:0]  adder_1_sub_2_io_s_delay_44;
  reg        [376:0]  adder_1_sub_2_io_s_delay_45;
  reg        [376:0]  adder_1_sub_2_io_s_delay_46;
  reg        [376:0]  adder_1_sub_2_io_s_delay_47;
  reg        [376:0]  adder_1_sub_2_io_s_delay_48;
  reg        [376:0]  adder_1_sub_2_io_s_delay_49;
  reg        [376:0]  adder_1_sub_2_io_s_delay_50;
  reg        [376:0]  adder_1_sub_2_io_s_delay_51;
  reg        [376:0]  adder_1_sub_2_io_s_delay_52;
  reg        [376:0]  adder_1_sub_2_io_s_delay_53;
  reg        [376:0]  adder_1_sub_2_io_s_delay_54;
  reg        [376:0]  adder_1_sub_2_io_s_delay_55;
  reg        [376:0]  adder_1_sub_2_io_s_delay_56;
  reg        [376:0]  adder_1_sub_2_io_s_delay_57;
  reg        [376:0]  adder_1_sub_2_io_s_delay_58;
  reg        [376:0]  adder_1_sub_2_io_s_delay_59;
  reg        [376:0]  adder_1_sub_2_io_s_delay_60;
  reg        [376:0]  adder_1_sub_2_io_s_delay_61;
  reg        [376:0]  adder_1_sub_2_io_s_delay_62;
  reg        [376:0]  adder_1_sub_2_io_s_delay_63;
  reg        [376:0]  adder_1_sub_2_io_s_delay_64;
  reg        [376:0]  adder_1_sub_2_io_s_delay_65;
  reg        [376:0]  adder_1_sub_2_io_s_delay_66;
  reg        [376:0]  adder_1_sub_2_io_s_delay_67;
  reg        [376:0]  adder_1_sub_2_io_s_delay_68;
  reg        [376:0]  adder_1_sub_2_io_s_delay_69;
  reg        [376:0]  adder_1_sub_2_io_s_delay_70;
  reg        [376:0]  adder_1_sub_2_io_s_delay_71;
  reg        [376:0]  adder_1_sub_2_io_s_delay_72;
  reg        [376:0]  adder_1_sub_2_io_s_delay_73;
  reg        [376:0]  adder_1_sub_2_io_s_delay_74;
  reg        [376:0]  adder_1_sub_2_io_s_delay_75;
  reg        [376:0]  R9;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_1;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_2;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_3;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_4;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_5;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_6;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_7;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_8;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_9;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_10;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_11;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_12;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_13;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_14;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_15;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_16;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_17;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_18;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_19;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_20;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_21;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_22;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_23;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_24;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_25;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_26;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_27;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_28;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_29;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_30;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_31;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_32;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_33;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_34;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_35;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_36;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_37;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_38;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_39;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_40;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_41;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_42;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_43;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_44;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_45;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_46;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_47;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_48;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_49;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_50;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_51;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_52;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_53;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_54;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_55;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_56;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_57;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_58;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_59;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_60;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_61;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_62;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_63;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_64;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_65;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_66;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_67;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_68;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_69;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_70;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_71;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_72;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_73;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_74;
  reg        [376:0]  adder_1_add_3_1_io_s_delay_75;
  reg        [376:0]  R12;

  KaratsubaMMUL_9 mul_0 (
    .io_a   (sub_0_io_s[376:0]), //i
    .io_b   (sub_1_io_s[376:0]), //i
    .io_p   (mul_0_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL_9 mul_1 (
    .io_a   (add_0_io_s[376:0]  ), //i
    .io_b   (add_1_1_io_s[376:0]), //i
    .io_p   (mul_1_io_p[376:0]  ), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  KaratsubaMMUL_9 mul_2 (
    .io_a   (io_a_T_delay_84[376:0]), //i
    .io_b   (cMul_io_p[376:0]      ), //i
    .io_p   (mul_2_io_p[376:0]     ), //o
    .clk    (clk                   ), //i
    .resetn (resetn                )  //i
  );
  KaratsubaMMUL_9 mul_3 (
    .io_a   (io_a_Z[376:0]    ), //i
    .io_b   (io_b_Z[376:0]    ), //i
    .io_p   (mul_3_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL_9 mul_4 (
    .io_a   (R9[376:0]        ), //i
    .io_b   (sub_3_io_s[376:0]), //i
    .io_p   (mul_4_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL_9 mul_5 (
    .io_a   (add_2_1_io_s[376:0]), //i
    .io_b   (R12[376:0]         ), //i
    .io_p   (mul_5_io_p[376:0]  ), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  KaratsubaMMUL_9 mul_6 (
    .io_a   (sub_3_io_s[376:0]  ), //i
    .io_b   (add_2_1_io_s[376:0]), //i
    .io_p   (mul_6_io_p[376:0]  ), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  KaratsubaMMUL_9 mul_7 (
    .io_a   (R9[376:0]        ), //i
    .io_b   (R12[376:0]       ), //i
    .io_p   (mul_7_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL_9 cMul (
    .io_a   (io_b_T[376:0]                                                                                       ), //i
    .io_b   (377'h196bab03169a4f2ca0b7670ae65fc7437786998c1a32d217f165b2fe0b32139735d947870e3d3e4e02c125684d6e016), //i
    .io_p   (cMul_io_p[376:0]                                                                                    ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  MADD_8 add_0 (
    .io_a   (io_a_Y[376:0]    ), //i
    .io_b   (io_a_X[376:0]    ), //i
    .io_s   (add_0_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_8 add_1_1 (
    .io_a   (io_b_Y[376:0]      ), //i
    .io_b   (io_b_X[376:0]      ), //i
    .io_s   (add_1_1_io_s[376:0]), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  MADD_8 add_2_1 (
    .io_a   (R8[376:0]          ), //i
    .io_b   (mul_2_io_p[376:0]  ), //i
    .io_s   (add_2_1_io_s[376:0]), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  MADD_8 add_3_1 (
    .io_a   (mul_1_io_p[376:0]  ), //i
    .io_b   (mul_0_io_p[376:0]  ), //i
    .io_s   (add_3_1_io_s[376:0]), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  MADD_12 sub_0 (
    .io_a   (io_a_Y[376:0]    ), //i
    .io_b   (io_a_X[376:0]    ), //i
    .io_s   (sub_0_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_12 sub_1 (
    .io_a   (io_b_Y[376:0]    ), //i
    .io_b   (io_b_X[376:0]    ), //i
    .io_s   (sub_1_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_12 sub_2 (
    .io_a   (mul_1_io_p[376:0]), //i
    .io_b   (mul_0_io_p[376:0]), //i
    .io_s   (sub_2_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_12 sub_3 (
    .io_a   (R8[376:0]        ), //i
    .io_b   (mul_2_io_p[376:0]), //i
    .io_s   (sub_3_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  FineReduction_1 reduction (
    .io_a   (reduction_io_a[377:0]), //i
    .io_r   (reduction_io_r[376:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign reduction_io_a = ({1'd0,mul_3_io_p} <<< 1);
  assign io_s_X = mul_4_io_p;
  assign io_s_Y = mul_5_io_p;
  assign io_s_Z = mul_6_io_p;
  assign io_s_T = mul_7_io_p;
  always @(posedge clk) begin
    io_a_T_delay_1 <= io_a_T;
    io_a_T_delay_2 <= io_a_T_delay_1;
    io_a_T_delay_3 <= io_a_T_delay_2;
    io_a_T_delay_4 <= io_a_T_delay_3;
    io_a_T_delay_5 <= io_a_T_delay_4;
    io_a_T_delay_6 <= io_a_T_delay_5;
    io_a_T_delay_7 <= io_a_T_delay_6;
    io_a_T_delay_8 <= io_a_T_delay_7;
    io_a_T_delay_9 <= io_a_T_delay_8;
    io_a_T_delay_10 <= io_a_T_delay_9;
    io_a_T_delay_11 <= io_a_T_delay_10;
    io_a_T_delay_12 <= io_a_T_delay_11;
    io_a_T_delay_13 <= io_a_T_delay_12;
    io_a_T_delay_14 <= io_a_T_delay_13;
    io_a_T_delay_15 <= io_a_T_delay_14;
    io_a_T_delay_16 <= io_a_T_delay_15;
    io_a_T_delay_17 <= io_a_T_delay_16;
    io_a_T_delay_18 <= io_a_T_delay_17;
    io_a_T_delay_19 <= io_a_T_delay_18;
    io_a_T_delay_20 <= io_a_T_delay_19;
    io_a_T_delay_21 <= io_a_T_delay_20;
    io_a_T_delay_22 <= io_a_T_delay_21;
    io_a_T_delay_23 <= io_a_T_delay_22;
    io_a_T_delay_24 <= io_a_T_delay_23;
    io_a_T_delay_25 <= io_a_T_delay_24;
    io_a_T_delay_26 <= io_a_T_delay_25;
    io_a_T_delay_27 <= io_a_T_delay_26;
    io_a_T_delay_28 <= io_a_T_delay_27;
    io_a_T_delay_29 <= io_a_T_delay_28;
    io_a_T_delay_30 <= io_a_T_delay_29;
    io_a_T_delay_31 <= io_a_T_delay_30;
    io_a_T_delay_32 <= io_a_T_delay_31;
    io_a_T_delay_33 <= io_a_T_delay_32;
    io_a_T_delay_34 <= io_a_T_delay_33;
    io_a_T_delay_35 <= io_a_T_delay_34;
    io_a_T_delay_36 <= io_a_T_delay_35;
    io_a_T_delay_37 <= io_a_T_delay_36;
    io_a_T_delay_38 <= io_a_T_delay_37;
    io_a_T_delay_39 <= io_a_T_delay_38;
    io_a_T_delay_40 <= io_a_T_delay_39;
    io_a_T_delay_41 <= io_a_T_delay_40;
    io_a_T_delay_42 <= io_a_T_delay_41;
    io_a_T_delay_43 <= io_a_T_delay_42;
    io_a_T_delay_44 <= io_a_T_delay_43;
    io_a_T_delay_45 <= io_a_T_delay_44;
    io_a_T_delay_46 <= io_a_T_delay_45;
    io_a_T_delay_47 <= io_a_T_delay_46;
    io_a_T_delay_48 <= io_a_T_delay_47;
    io_a_T_delay_49 <= io_a_T_delay_48;
    io_a_T_delay_50 <= io_a_T_delay_49;
    io_a_T_delay_51 <= io_a_T_delay_50;
    io_a_T_delay_52 <= io_a_T_delay_51;
    io_a_T_delay_53 <= io_a_T_delay_52;
    io_a_T_delay_54 <= io_a_T_delay_53;
    io_a_T_delay_55 <= io_a_T_delay_54;
    io_a_T_delay_56 <= io_a_T_delay_55;
    io_a_T_delay_57 <= io_a_T_delay_56;
    io_a_T_delay_58 <= io_a_T_delay_57;
    io_a_T_delay_59 <= io_a_T_delay_58;
    io_a_T_delay_60 <= io_a_T_delay_59;
    io_a_T_delay_61 <= io_a_T_delay_60;
    io_a_T_delay_62 <= io_a_T_delay_61;
    io_a_T_delay_63 <= io_a_T_delay_62;
    io_a_T_delay_64 <= io_a_T_delay_63;
    io_a_T_delay_65 <= io_a_T_delay_64;
    io_a_T_delay_66 <= io_a_T_delay_65;
    io_a_T_delay_67 <= io_a_T_delay_66;
    io_a_T_delay_68 <= io_a_T_delay_67;
    io_a_T_delay_69 <= io_a_T_delay_68;
    io_a_T_delay_70 <= io_a_T_delay_69;
    io_a_T_delay_71 <= io_a_T_delay_70;
    io_a_T_delay_72 <= io_a_T_delay_71;
    io_a_T_delay_73 <= io_a_T_delay_72;
    io_a_T_delay_74 <= io_a_T_delay_73;
    io_a_T_delay_75 <= io_a_T_delay_74;
    io_a_T_delay_76 <= io_a_T_delay_75;
    io_a_T_delay_77 <= io_a_T_delay_76;
    io_a_T_delay_78 <= io_a_T_delay_77;
    io_a_T_delay_79 <= io_a_T_delay_78;
    io_a_T_delay_80 <= io_a_T_delay_79;
    io_a_T_delay_81 <= io_a_T_delay_80;
    io_a_T_delay_82 <= io_a_T_delay_81;
    io_a_T_delay_83 <= io_a_T_delay_82;
    io_a_T_delay_84 <= io_a_T_delay_83;
    adder_1_reduction_io_r_delay_1 <= reduction_io_r;
    adder_1_reduction_io_r_delay_2 <= adder_1_reduction_io_r_delay_1;
    adder_1_reduction_io_r_delay_3 <= adder_1_reduction_io_r_delay_2;
    adder_1_reduction_io_r_delay_4 <= adder_1_reduction_io_r_delay_3;
    adder_1_reduction_io_r_delay_5 <= adder_1_reduction_io_r_delay_4;
    adder_1_reduction_io_r_delay_6 <= adder_1_reduction_io_r_delay_5;
    adder_1_reduction_io_r_delay_7 <= adder_1_reduction_io_r_delay_6;
    adder_1_reduction_io_r_delay_8 <= adder_1_reduction_io_r_delay_7;
    adder_1_reduction_io_r_delay_9 <= adder_1_reduction_io_r_delay_8;
    adder_1_reduction_io_r_delay_10 <= adder_1_reduction_io_r_delay_9;
    adder_1_reduction_io_r_delay_11 <= adder_1_reduction_io_r_delay_10;
    adder_1_reduction_io_r_delay_12 <= adder_1_reduction_io_r_delay_11;
    adder_1_reduction_io_r_delay_13 <= adder_1_reduction_io_r_delay_12;
    adder_1_reduction_io_r_delay_14 <= adder_1_reduction_io_r_delay_13;
    adder_1_reduction_io_r_delay_15 <= adder_1_reduction_io_r_delay_14;
    adder_1_reduction_io_r_delay_16 <= adder_1_reduction_io_r_delay_15;
    adder_1_reduction_io_r_delay_17 <= adder_1_reduction_io_r_delay_16;
    adder_1_reduction_io_r_delay_18 <= adder_1_reduction_io_r_delay_17;
    adder_1_reduction_io_r_delay_19 <= adder_1_reduction_io_r_delay_18;
    adder_1_reduction_io_r_delay_20 <= adder_1_reduction_io_r_delay_19;
    adder_1_reduction_io_r_delay_21 <= adder_1_reduction_io_r_delay_20;
    adder_1_reduction_io_r_delay_22 <= adder_1_reduction_io_r_delay_21;
    adder_1_reduction_io_r_delay_23 <= adder_1_reduction_io_r_delay_22;
    adder_1_reduction_io_r_delay_24 <= adder_1_reduction_io_r_delay_23;
    adder_1_reduction_io_r_delay_25 <= adder_1_reduction_io_r_delay_24;
    adder_1_reduction_io_r_delay_26 <= adder_1_reduction_io_r_delay_25;
    adder_1_reduction_io_r_delay_27 <= adder_1_reduction_io_r_delay_26;
    adder_1_reduction_io_r_delay_28 <= adder_1_reduction_io_r_delay_27;
    adder_1_reduction_io_r_delay_29 <= adder_1_reduction_io_r_delay_28;
    adder_1_reduction_io_r_delay_30 <= adder_1_reduction_io_r_delay_29;
    adder_1_reduction_io_r_delay_31 <= adder_1_reduction_io_r_delay_30;
    adder_1_reduction_io_r_delay_32 <= adder_1_reduction_io_r_delay_31;
    adder_1_reduction_io_r_delay_33 <= adder_1_reduction_io_r_delay_32;
    adder_1_reduction_io_r_delay_34 <= adder_1_reduction_io_r_delay_33;
    adder_1_reduction_io_r_delay_35 <= adder_1_reduction_io_r_delay_34;
    adder_1_reduction_io_r_delay_36 <= adder_1_reduction_io_r_delay_35;
    adder_1_reduction_io_r_delay_37 <= adder_1_reduction_io_r_delay_36;
    adder_1_reduction_io_r_delay_38 <= adder_1_reduction_io_r_delay_37;
    adder_1_reduction_io_r_delay_39 <= adder_1_reduction_io_r_delay_38;
    adder_1_reduction_io_r_delay_40 <= adder_1_reduction_io_r_delay_39;
    adder_1_reduction_io_r_delay_41 <= adder_1_reduction_io_r_delay_40;
    adder_1_reduction_io_r_delay_42 <= adder_1_reduction_io_r_delay_41;
    adder_1_reduction_io_r_delay_43 <= adder_1_reduction_io_r_delay_42;
    adder_1_reduction_io_r_delay_44 <= adder_1_reduction_io_r_delay_43;
    adder_1_reduction_io_r_delay_45 <= adder_1_reduction_io_r_delay_44;
    adder_1_reduction_io_r_delay_46 <= adder_1_reduction_io_r_delay_45;
    adder_1_reduction_io_r_delay_47 <= adder_1_reduction_io_r_delay_46;
    adder_1_reduction_io_r_delay_48 <= adder_1_reduction_io_r_delay_47;
    adder_1_reduction_io_r_delay_49 <= adder_1_reduction_io_r_delay_48;
    adder_1_reduction_io_r_delay_50 <= adder_1_reduction_io_r_delay_49;
    adder_1_reduction_io_r_delay_51 <= adder_1_reduction_io_r_delay_50;
    adder_1_reduction_io_r_delay_52 <= adder_1_reduction_io_r_delay_51;
    adder_1_reduction_io_r_delay_53 <= adder_1_reduction_io_r_delay_52;
    adder_1_reduction_io_r_delay_54 <= adder_1_reduction_io_r_delay_53;
    adder_1_reduction_io_r_delay_55 <= adder_1_reduction_io_r_delay_54;
    adder_1_reduction_io_r_delay_56 <= adder_1_reduction_io_r_delay_55;
    adder_1_reduction_io_r_delay_57 <= adder_1_reduction_io_r_delay_56;
    adder_1_reduction_io_r_delay_58 <= adder_1_reduction_io_r_delay_57;
    adder_1_reduction_io_r_delay_59 <= adder_1_reduction_io_r_delay_58;
    adder_1_reduction_io_r_delay_60 <= adder_1_reduction_io_r_delay_59;
    adder_1_reduction_io_r_delay_61 <= adder_1_reduction_io_r_delay_60;
    adder_1_reduction_io_r_delay_62 <= adder_1_reduction_io_r_delay_61;
    adder_1_reduction_io_r_delay_63 <= adder_1_reduction_io_r_delay_62;
    adder_1_reduction_io_r_delay_64 <= adder_1_reduction_io_r_delay_63;
    adder_1_reduction_io_r_delay_65 <= adder_1_reduction_io_r_delay_64;
    adder_1_reduction_io_r_delay_66 <= adder_1_reduction_io_r_delay_65;
    adder_1_reduction_io_r_delay_67 <= adder_1_reduction_io_r_delay_66;
    adder_1_reduction_io_r_delay_68 <= adder_1_reduction_io_r_delay_67;
    adder_1_reduction_io_r_delay_69 <= adder_1_reduction_io_r_delay_68;
    adder_1_reduction_io_r_delay_70 <= adder_1_reduction_io_r_delay_69;
    adder_1_reduction_io_r_delay_71 <= adder_1_reduction_io_r_delay_70;
    adder_1_reduction_io_r_delay_72 <= adder_1_reduction_io_r_delay_71;
    adder_1_reduction_io_r_delay_73 <= adder_1_reduction_io_r_delay_72;
    adder_1_reduction_io_r_delay_74 <= adder_1_reduction_io_r_delay_73;
    adder_1_reduction_io_r_delay_75 <= adder_1_reduction_io_r_delay_74;
    adder_1_reduction_io_r_delay_76 <= adder_1_reduction_io_r_delay_75;
    R8 <= adder_1_reduction_io_r_delay_76;
    adder_1_sub_2_io_s_delay_1 <= sub_2_io_s;
    adder_1_sub_2_io_s_delay_2 <= adder_1_sub_2_io_s_delay_1;
    adder_1_sub_2_io_s_delay_3 <= adder_1_sub_2_io_s_delay_2;
    adder_1_sub_2_io_s_delay_4 <= adder_1_sub_2_io_s_delay_3;
    adder_1_sub_2_io_s_delay_5 <= adder_1_sub_2_io_s_delay_4;
    adder_1_sub_2_io_s_delay_6 <= adder_1_sub_2_io_s_delay_5;
    adder_1_sub_2_io_s_delay_7 <= adder_1_sub_2_io_s_delay_6;
    adder_1_sub_2_io_s_delay_8 <= adder_1_sub_2_io_s_delay_7;
    adder_1_sub_2_io_s_delay_9 <= adder_1_sub_2_io_s_delay_8;
    adder_1_sub_2_io_s_delay_10 <= adder_1_sub_2_io_s_delay_9;
    adder_1_sub_2_io_s_delay_11 <= adder_1_sub_2_io_s_delay_10;
    adder_1_sub_2_io_s_delay_12 <= adder_1_sub_2_io_s_delay_11;
    adder_1_sub_2_io_s_delay_13 <= adder_1_sub_2_io_s_delay_12;
    adder_1_sub_2_io_s_delay_14 <= adder_1_sub_2_io_s_delay_13;
    adder_1_sub_2_io_s_delay_15 <= adder_1_sub_2_io_s_delay_14;
    adder_1_sub_2_io_s_delay_16 <= adder_1_sub_2_io_s_delay_15;
    adder_1_sub_2_io_s_delay_17 <= adder_1_sub_2_io_s_delay_16;
    adder_1_sub_2_io_s_delay_18 <= adder_1_sub_2_io_s_delay_17;
    adder_1_sub_2_io_s_delay_19 <= adder_1_sub_2_io_s_delay_18;
    adder_1_sub_2_io_s_delay_20 <= adder_1_sub_2_io_s_delay_19;
    adder_1_sub_2_io_s_delay_21 <= adder_1_sub_2_io_s_delay_20;
    adder_1_sub_2_io_s_delay_22 <= adder_1_sub_2_io_s_delay_21;
    adder_1_sub_2_io_s_delay_23 <= adder_1_sub_2_io_s_delay_22;
    adder_1_sub_2_io_s_delay_24 <= adder_1_sub_2_io_s_delay_23;
    adder_1_sub_2_io_s_delay_25 <= adder_1_sub_2_io_s_delay_24;
    adder_1_sub_2_io_s_delay_26 <= adder_1_sub_2_io_s_delay_25;
    adder_1_sub_2_io_s_delay_27 <= adder_1_sub_2_io_s_delay_26;
    adder_1_sub_2_io_s_delay_28 <= adder_1_sub_2_io_s_delay_27;
    adder_1_sub_2_io_s_delay_29 <= adder_1_sub_2_io_s_delay_28;
    adder_1_sub_2_io_s_delay_30 <= adder_1_sub_2_io_s_delay_29;
    adder_1_sub_2_io_s_delay_31 <= adder_1_sub_2_io_s_delay_30;
    adder_1_sub_2_io_s_delay_32 <= adder_1_sub_2_io_s_delay_31;
    adder_1_sub_2_io_s_delay_33 <= adder_1_sub_2_io_s_delay_32;
    adder_1_sub_2_io_s_delay_34 <= adder_1_sub_2_io_s_delay_33;
    adder_1_sub_2_io_s_delay_35 <= adder_1_sub_2_io_s_delay_34;
    adder_1_sub_2_io_s_delay_36 <= adder_1_sub_2_io_s_delay_35;
    adder_1_sub_2_io_s_delay_37 <= adder_1_sub_2_io_s_delay_36;
    adder_1_sub_2_io_s_delay_38 <= adder_1_sub_2_io_s_delay_37;
    adder_1_sub_2_io_s_delay_39 <= adder_1_sub_2_io_s_delay_38;
    adder_1_sub_2_io_s_delay_40 <= adder_1_sub_2_io_s_delay_39;
    adder_1_sub_2_io_s_delay_41 <= adder_1_sub_2_io_s_delay_40;
    adder_1_sub_2_io_s_delay_42 <= adder_1_sub_2_io_s_delay_41;
    adder_1_sub_2_io_s_delay_43 <= adder_1_sub_2_io_s_delay_42;
    adder_1_sub_2_io_s_delay_44 <= adder_1_sub_2_io_s_delay_43;
    adder_1_sub_2_io_s_delay_45 <= adder_1_sub_2_io_s_delay_44;
    adder_1_sub_2_io_s_delay_46 <= adder_1_sub_2_io_s_delay_45;
    adder_1_sub_2_io_s_delay_47 <= adder_1_sub_2_io_s_delay_46;
    adder_1_sub_2_io_s_delay_48 <= adder_1_sub_2_io_s_delay_47;
    adder_1_sub_2_io_s_delay_49 <= adder_1_sub_2_io_s_delay_48;
    adder_1_sub_2_io_s_delay_50 <= adder_1_sub_2_io_s_delay_49;
    adder_1_sub_2_io_s_delay_51 <= adder_1_sub_2_io_s_delay_50;
    adder_1_sub_2_io_s_delay_52 <= adder_1_sub_2_io_s_delay_51;
    adder_1_sub_2_io_s_delay_53 <= adder_1_sub_2_io_s_delay_52;
    adder_1_sub_2_io_s_delay_54 <= adder_1_sub_2_io_s_delay_53;
    adder_1_sub_2_io_s_delay_55 <= adder_1_sub_2_io_s_delay_54;
    adder_1_sub_2_io_s_delay_56 <= adder_1_sub_2_io_s_delay_55;
    adder_1_sub_2_io_s_delay_57 <= adder_1_sub_2_io_s_delay_56;
    adder_1_sub_2_io_s_delay_58 <= adder_1_sub_2_io_s_delay_57;
    adder_1_sub_2_io_s_delay_59 <= adder_1_sub_2_io_s_delay_58;
    adder_1_sub_2_io_s_delay_60 <= adder_1_sub_2_io_s_delay_59;
    adder_1_sub_2_io_s_delay_61 <= adder_1_sub_2_io_s_delay_60;
    adder_1_sub_2_io_s_delay_62 <= adder_1_sub_2_io_s_delay_61;
    adder_1_sub_2_io_s_delay_63 <= adder_1_sub_2_io_s_delay_62;
    adder_1_sub_2_io_s_delay_64 <= adder_1_sub_2_io_s_delay_63;
    adder_1_sub_2_io_s_delay_65 <= adder_1_sub_2_io_s_delay_64;
    adder_1_sub_2_io_s_delay_66 <= adder_1_sub_2_io_s_delay_65;
    adder_1_sub_2_io_s_delay_67 <= adder_1_sub_2_io_s_delay_66;
    adder_1_sub_2_io_s_delay_68 <= adder_1_sub_2_io_s_delay_67;
    adder_1_sub_2_io_s_delay_69 <= adder_1_sub_2_io_s_delay_68;
    adder_1_sub_2_io_s_delay_70 <= adder_1_sub_2_io_s_delay_69;
    adder_1_sub_2_io_s_delay_71 <= adder_1_sub_2_io_s_delay_70;
    adder_1_sub_2_io_s_delay_72 <= adder_1_sub_2_io_s_delay_71;
    adder_1_sub_2_io_s_delay_73 <= adder_1_sub_2_io_s_delay_72;
    adder_1_sub_2_io_s_delay_74 <= adder_1_sub_2_io_s_delay_73;
    adder_1_sub_2_io_s_delay_75 <= adder_1_sub_2_io_s_delay_74;
    R9 <= adder_1_sub_2_io_s_delay_75;
    adder_1_add_3_1_io_s_delay_1 <= add_3_1_io_s;
    adder_1_add_3_1_io_s_delay_2 <= adder_1_add_3_1_io_s_delay_1;
    adder_1_add_3_1_io_s_delay_3 <= adder_1_add_3_1_io_s_delay_2;
    adder_1_add_3_1_io_s_delay_4 <= adder_1_add_3_1_io_s_delay_3;
    adder_1_add_3_1_io_s_delay_5 <= adder_1_add_3_1_io_s_delay_4;
    adder_1_add_3_1_io_s_delay_6 <= adder_1_add_3_1_io_s_delay_5;
    adder_1_add_3_1_io_s_delay_7 <= adder_1_add_3_1_io_s_delay_6;
    adder_1_add_3_1_io_s_delay_8 <= adder_1_add_3_1_io_s_delay_7;
    adder_1_add_3_1_io_s_delay_9 <= adder_1_add_3_1_io_s_delay_8;
    adder_1_add_3_1_io_s_delay_10 <= adder_1_add_3_1_io_s_delay_9;
    adder_1_add_3_1_io_s_delay_11 <= adder_1_add_3_1_io_s_delay_10;
    adder_1_add_3_1_io_s_delay_12 <= adder_1_add_3_1_io_s_delay_11;
    adder_1_add_3_1_io_s_delay_13 <= adder_1_add_3_1_io_s_delay_12;
    adder_1_add_3_1_io_s_delay_14 <= adder_1_add_3_1_io_s_delay_13;
    adder_1_add_3_1_io_s_delay_15 <= adder_1_add_3_1_io_s_delay_14;
    adder_1_add_3_1_io_s_delay_16 <= adder_1_add_3_1_io_s_delay_15;
    adder_1_add_3_1_io_s_delay_17 <= adder_1_add_3_1_io_s_delay_16;
    adder_1_add_3_1_io_s_delay_18 <= adder_1_add_3_1_io_s_delay_17;
    adder_1_add_3_1_io_s_delay_19 <= adder_1_add_3_1_io_s_delay_18;
    adder_1_add_3_1_io_s_delay_20 <= adder_1_add_3_1_io_s_delay_19;
    adder_1_add_3_1_io_s_delay_21 <= adder_1_add_3_1_io_s_delay_20;
    adder_1_add_3_1_io_s_delay_22 <= adder_1_add_3_1_io_s_delay_21;
    adder_1_add_3_1_io_s_delay_23 <= adder_1_add_3_1_io_s_delay_22;
    adder_1_add_3_1_io_s_delay_24 <= adder_1_add_3_1_io_s_delay_23;
    adder_1_add_3_1_io_s_delay_25 <= adder_1_add_3_1_io_s_delay_24;
    adder_1_add_3_1_io_s_delay_26 <= adder_1_add_3_1_io_s_delay_25;
    adder_1_add_3_1_io_s_delay_27 <= adder_1_add_3_1_io_s_delay_26;
    adder_1_add_3_1_io_s_delay_28 <= adder_1_add_3_1_io_s_delay_27;
    adder_1_add_3_1_io_s_delay_29 <= adder_1_add_3_1_io_s_delay_28;
    adder_1_add_3_1_io_s_delay_30 <= adder_1_add_3_1_io_s_delay_29;
    adder_1_add_3_1_io_s_delay_31 <= adder_1_add_3_1_io_s_delay_30;
    adder_1_add_3_1_io_s_delay_32 <= adder_1_add_3_1_io_s_delay_31;
    adder_1_add_3_1_io_s_delay_33 <= adder_1_add_3_1_io_s_delay_32;
    adder_1_add_3_1_io_s_delay_34 <= adder_1_add_3_1_io_s_delay_33;
    adder_1_add_3_1_io_s_delay_35 <= adder_1_add_3_1_io_s_delay_34;
    adder_1_add_3_1_io_s_delay_36 <= adder_1_add_3_1_io_s_delay_35;
    adder_1_add_3_1_io_s_delay_37 <= adder_1_add_3_1_io_s_delay_36;
    adder_1_add_3_1_io_s_delay_38 <= adder_1_add_3_1_io_s_delay_37;
    adder_1_add_3_1_io_s_delay_39 <= adder_1_add_3_1_io_s_delay_38;
    adder_1_add_3_1_io_s_delay_40 <= adder_1_add_3_1_io_s_delay_39;
    adder_1_add_3_1_io_s_delay_41 <= adder_1_add_3_1_io_s_delay_40;
    adder_1_add_3_1_io_s_delay_42 <= adder_1_add_3_1_io_s_delay_41;
    adder_1_add_3_1_io_s_delay_43 <= adder_1_add_3_1_io_s_delay_42;
    adder_1_add_3_1_io_s_delay_44 <= adder_1_add_3_1_io_s_delay_43;
    adder_1_add_3_1_io_s_delay_45 <= adder_1_add_3_1_io_s_delay_44;
    adder_1_add_3_1_io_s_delay_46 <= adder_1_add_3_1_io_s_delay_45;
    adder_1_add_3_1_io_s_delay_47 <= adder_1_add_3_1_io_s_delay_46;
    adder_1_add_3_1_io_s_delay_48 <= adder_1_add_3_1_io_s_delay_47;
    adder_1_add_3_1_io_s_delay_49 <= adder_1_add_3_1_io_s_delay_48;
    adder_1_add_3_1_io_s_delay_50 <= adder_1_add_3_1_io_s_delay_49;
    adder_1_add_3_1_io_s_delay_51 <= adder_1_add_3_1_io_s_delay_50;
    adder_1_add_3_1_io_s_delay_52 <= adder_1_add_3_1_io_s_delay_51;
    adder_1_add_3_1_io_s_delay_53 <= adder_1_add_3_1_io_s_delay_52;
    adder_1_add_3_1_io_s_delay_54 <= adder_1_add_3_1_io_s_delay_53;
    adder_1_add_3_1_io_s_delay_55 <= adder_1_add_3_1_io_s_delay_54;
    adder_1_add_3_1_io_s_delay_56 <= adder_1_add_3_1_io_s_delay_55;
    adder_1_add_3_1_io_s_delay_57 <= adder_1_add_3_1_io_s_delay_56;
    adder_1_add_3_1_io_s_delay_58 <= adder_1_add_3_1_io_s_delay_57;
    adder_1_add_3_1_io_s_delay_59 <= adder_1_add_3_1_io_s_delay_58;
    adder_1_add_3_1_io_s_delay_60 <= adder_1_add_3_1_io_s_delay_59;
    adder_1_add_3_1_io_s_delay_61 <= adder_1_add_3_1_io_s_delay_60;
    adder_1_add_3_1_io_s_delay_62 <= adder_1_add_3_1_io_s_delay_61;
    adder_1_add_3_1_io_s_delay_63 <= adder_1_add_3_1_io_s_delay_62;
    adder_1_add_3_1_io_s_delay_64 <= adder_1_add_3_1_io_s_delay_63;
    adder_1_add_3_1_io_s_delay_65 <= adder_1_add_3_1_io_s_delay_64;
    adder_1_add_3_1_io_s_delay_66 <= adder_1_add_3_1_io_s_delay_65;
    adder_1_add_3_1_io_s_delay_67 <= adder_1_add_3_1_io_s_delay_66;
    adder_1_add_3_1_io_s_delay_68 <= adder_1_add_3_1_io_s_delay_67;
    adder_1_add_3_1_io_s_delay_69 <= adder_1_add_3_1_io_s_delay_68;
    adder_1_add_3_1_io_s_delay_70 <= adder_1_add_3_1_io_s_delay_69;
    adder_1_add_3_1_io_s_delay_71 <= adder_1_add_3_1_io_s_delay_70;
    adder_1_add_3_1_io_s_delay_72 <= adder_1_add_3_1_io_s_delay_71;
    adder_1_add_3_1_io_s_delay_73 <= adder_1_add_3_1_io_s_delay_72;
    adder_1_add_3_1_io_s_delay_74 <= adder_1_add_3_1_io_s_delay_73;
    adder_1_add_3_1_io_s_delay_75 <= adder_1_add_3_1_io_s_delay_74;
    R12 <= adder_1_add_3_1_io_s_delay_75;
  end


endmodule

module PAdd (
  input      [376:0]  io_a_X,
  input      [376:0]  io_a_Y,
  input      [376:0]  io_a_Z,
  input      [376:0]  io_a_T,
  input      [376:0]  io_b_X,
  input      [376:0]  io_b_Y,
  input      [376:0]  io_b_Z,
  input      [376:0]  io_b_T,
  output     [376:0]  io_s_X,
  output     [376:0]  io_s_Y,
  output     [376:0]  io_s_Z,
  output     [376:0]  io_s_T,
  input               clk,
  input               resetn
);

  wire       [377:0]  reduction_io_a;
  wire       [376:0]  mul_0_io_p;
  wire       [376:0]  mul_1_io_p;
  wire       [376:0]  mul_2_io_p;
  wire       [376:0]  mul_3_io_p;
  wire       [376:0]  mul_4_io_p;
  wire       [376:0]  mul_5_io_p;
  wire       [376:0]  mul_6_io_p;
  wire       [376:0]  mul_7_io_p;
  wire       [376:0]  cMul_io_p;
  wire       [376:0]  add_0_io_s;
  wire       [376:0]  add_1_1_io_s;
  wire       [376:0]  add_2_1_io_s;
  wire       [376:0]  add_3_1_io_s;
  wire       [376:0]  sub_0_io_s;
  wire       [376:0]  sub_1_io_s;
  wire       [376:0]  sub_2_io_s;
  wire       [376:0]  sub_3_io_s;
  wire       [376:0]  reduction_io_r;
  reg        [376:0]  io_a_T_delay_1;
  reg        [376:0]  io_a_T_delay_2;
  reg        [376:0]  io_a_T_delay_3;
  reg        [376:0]  io_a_T_delay_4;
  reg        [376:0]  io_a_T_delay_5;
  reg        [376:0]  io_a_T_delay_6;
  reg        [376:0]  io_a_T_delay_7;
  reg        [376:0]  io_a_T_delay_8;
  reg        [376:0]  io_a_T_delay_9;
  reg        [376:0]  io_a_T_delay_10;
  reg        [376:0]  io_a_T_delay_11;
  reg        [376:0]  io_a_T_delay_12;
  reg        [376:0]  io_a_T_delay_13;
  reg        [376:0]  io_a_T_delay_14;
  reg        [376:0]  io_a_T_delay_15;
  reg        [376:0]  io_a_T_delay_16;
  reg        [376:0]  io_a_T_delay_17;
  reg        [376:0]  io_a_T_delay_18;
  reg        [376:0]  io_a_T_delay_19;
  reg        [376:0]  io_a_T_delay_20;
  reg        [376:0]  io_a_T_delay_21;
  reg        [376:0]  io_a_T_delay_22;
  reg        [376:0]  io_a_T_delay_23;
  reg        [376:0]  io_a_T_delay_24;
  reg        [376:0]  io_a_T_delay_25;
  reg        [376:0]  io_a_T_delay_26;
  reg        [376:0]  io_a_T_delay_27;
  reg        [376:0]  io_a_T_delay_28;
  reg        [376:0]  io_a_T_delay_29;
  reg        [376:0]  io_a_T_delay_30;
  reg        [376:0]  io_a_T_delay_31;
  reg        [376:0]  io_a_T_delay_32;
  reg        [376:0]  io_a_T_delay_33;
  reg        [376:0]  io_a_T_delay_34;
  reg        [376:0]  io_a_T_delay_35;
  reg        [376:0]  io_a_T_delay_36;
  reg        [376:0]  io_a_T_delay_37;
  reg        [376:0]  io_a_T_delay_38;
  reg        [376:0]  io_a_T_delay_39;
  reg        [376:0]  io_a_T_delay_40;
  reg        [376:0]  io_a_T_delay_41;
  reg        [376:0]  io_a_T_delay_42;
  reg        [376:0]  io_a_T_delay_43;
  reg        [376:0]  io_a_T_delay_44;
  reg        [376:0]  io_a_T_delay_45;
  reg        [376:0]  io_a_T_delay_46;
  reg        [376:0]  io_a_T_delay_47;
  reg        [376:0]  io_a_T_delay_48;
  reg        [376:0]  io_a_T_delay_49;
  reg        [376:0]  io_a_T_delay_50;
  reg        [376:0]  io_a_T_delay_51;
  reg        [376:0]  io_a_T_delay_52;
  reg        [376:0]  io_a_T_delay_53;
  reg        [376:0]  io_a_T_delay_54;
  reg        [376:0]  io_a_T_delay_55;
  reg        [376:0]  io_a_T_delay_56;
  reg        [376:0]  io_a_T_delay_57;
  reg        [376:0]  io_a_T_delay_58;
  reg        [376:0]  io_a_T_delay_59;
  reg        [376:0]  io_a_T_delay_60;
  reg        [376:0]  io_a_T_delay_61;
  reg        [376:0]  io_a_T_delay_62;
  reg        [376:0]  io_a_T_delay_63;
  reg        [376:0]  io_a_T_delay_64;
  reg        [376:0]  io_a_T_delay_65;
  reg        [376:0]  io_a_T_delay_66;
  reg        [376:0]  io_a_T_delay_67;
  reg        [376:0]  io_a_T_delay_68;
  reg        [376:0]  io_a_T_delay_69;
  reg        [376:0]  io_a_T_delay_70;
  reg        [376:0]  io_a_T_delay_71;
  reg        [376:0]  io_a_T_delay_72;
  reg        [376:0]  io_a_T_delay_73;
  reg        [376:0]  io_a_T_delay_74;
  reg        [376:0]  io_a_T_delay_75;
  reg        [376:0]  io_a_T_delay_76;
  reg        [376:0]  io_a_T_delay_77;
  reg        [376:0]  io_a_T_delay_78;
  reg        [376:0]  io_a_T_delay_79;
  reg        [376:0]  io_a_T_delay_80;
  reg        [376:0]  io_a_T_delay_81;
  reg        [376:0]  io_a_T_delay_82;
  reg        [376:0]  io_a_T_delay_83;
  reg        [376:0]  io_a_T_delay_84;
  reg        [376:0]  adder_0_reduction_io_r_delay_1;
  reg        [376:0]  adder_0_reduction_io_r_delay_2;
  reg        [376:0]  adder_0_reduction_io_r_delay_3;
  reg        [376:0]  adder_0_reduction_io_r_delay_4;
  reg        [376:0]  adder_0_reduction_io_r_delay_5;
  reg        [376:0]  adder_0_reduction_io_r_delay_6;
  reg        [376:0]  adder_0_reduction_io_r_delay_7;
  reg        [376:0]  adder_0_reduction_io_r_delay_8;
  reg        [376:0]  adder_0_reduction_io_r_delay_9;
  reg        [376:0]  adder_0_reduction_io_r_delay_10;
  reg        [376:0]  adder_0_reduction_io_r_delay_11;
  reg        [376:0]  adder_0_reduction_io_r_delay_12;
  reg        [376:0]  adder_0_reduction_io_r_delay_13;
  reg        [376:0]  adder_0_reduction_io_r_delay_14;
  reg        [376:0]  adder_0_reduction_io_r_delay_15;
  reg        [376:0]  adder_0_reduction_io_r_delay_16;
  reg        [376:0]  adder_0_reduction_io_r_delay_17;
  reg        [376:0]  adder_0_reduction_io_r_delay_18;
  reg        [376:0]  adder_0_reduction_io_r_delay_19;
  reg        [376:0]  adder_0_reduction_io_r_delay_20;
  reg        [376:0]  adder_0_reduction_io_r_delay_21;
  reg        [376:0]  adder_0_reduction_io_r_delay_22;
  reg        [376:0]  adder_0_reduction_io_r_delay_23;
  reg        [376:0]  adder_0_reduction_io_r_delay_24;
  reg        [376:0]  adder_0_reduction_io_r_delay_25;
  reg        [376:0]  adder_0_reduction_io_r_delay_26;
  reg        [376:0]  adder_0_reduction_io_r_delay_27;
  reg        [376:0]  adder_0_reduction_io_r_delay_28;
  reg        [376:0]  adder_0_reduction_io_r_delay_29;
  reg        [376:0]  adder_0_reduction_io_r_delay_30;
  reg        [376:0]  adder_0_reduction_io_r_delay_31;
  reg        [376:0]  adder_0_reduction_io_r_delay_32;
  reg        [376:0]  adder_0_reduction_io_r_delay_33;
  reg        [376:0]  adder_0_reduction_io_r_delay_34;
  reg        [376:0]  adder_0_reduction_io_r_delay_35;
  reg        [376:0]  adder_0_reduction_io_r_delay_36;
  reg        [376:0]  adder_0_reduction_io_r_delay_37;
  reg        [376:0]  adder_0_reduction_io_r_delay_38;
  reg        [376:0]  adder_0_reduction_io_r_delay_39;
  reg        [376:0]  adder_0_reduction_io_r_delay_40;
  reg        [376:0]  adder_0_reduction_io_r_delay_41;
  reg        [376:0]  adder_0_reduction_io_r_delay_42;
  reg        [376:0]  adder_0_reduction_io_r_delay_43;
  reg        [376:0]  adder_0_reduction_io_r_delay_44;
  reg        [376:0]  adder_0_reduction_io_r_delay_45;
  reg        [376:0]  adder_0_reduction_io_r_delay_46;
  reg        [376:0]  adder_0_reduction_io_r_delay_47;
  reg        [376:0]  adder_0_reduction_io_r_delay_48;
  reg        [376:0]  adder_0_reduction_io_r_delay_49;
  reg        [376:0]  adder_0_reduction_io_r_delay_50;
  reg        [376:0]  adder_0_reduction_io_r_delay_51;
  reg        [376:0]  adder_0_reduction_io_r_delay_52;
  reg        [376:0]  adder_0_reduction_io_r_delay_53;
  reg        [376:0]  adder_0_reduction_io_r_delay_54;
  reg        [376:0]  adder_0_reduction_io_r_delay_55;
  reg        [376:0]  adder_0_reduction_io_r_delay_56;
  reg        [376:0]  adder_0_reduction_io_r_delay_57;
  reg        [376:0]  adder_0_reduction_io_r_delay_58;
  reg        [376:0]  adder_0_reduction_io_r_delay_59;
  reg        [376:0]  adder_0_reduction_io_r_delay_60;
  reg        [376:0]  adder_0_reduction_io_r_delay_61;
  reg        [376:0]  adder_0_reduction_io_r_delay_62;
  reg        [376:0]  adder_0_reduction_io_r_delay_63;
  reg        [376:0]  adder_0_reduction_io_r_delay_64;
  reg        [376:0]  adder_0_reduction_io_r_delay_65;
  reg        [376:0]  adder_0_reduction_io_r_delay_66;
  reg        [376:0]  adder_0_reduction_io_r_delay_67;
  reg        [376:0]  adder_0_reduction_io_r_delay_68;
  reg        [376:0]  adder_0_reduction_io_r_delay_69;
  reg        [376:0]  adder_0_reduction_io_r_delay_70;
  reg        [376:0]  adder_0_reduction_io_r_delay_71;
  reg        [376:0]  adder_0_reduction_io_r_delay_72;
  reg        [376:0]  adder_0_reduction_io_r_delay_73;
  reg        [376:0]  adder_0_reduction_io_r_delay_74;
  reg        [376:0]  adder_0_reduction_io_r_delay_75;
  reg        [376:0]  adder_0_reduction_io_r_delay_76;
  reg        [376:0]  R8;
  reg        [376:0]  adder_0_sub_2_io_s_delay_1;
  reg        [376:0]  adder_0_sub_2_io_s_delay_2;
  reg        [376:0]  adder_0_sub_2_io_s_delay_3;
  reg        [376:0]  adder_0_sub_2_io_s_delay_4;
  reg        [376:0]  adder_0_sub_2_io_s_delay_5;
  reg        [376:0]  adder_0_sub_2_io_s_delay_6;
  reg        [376:0]  adder_0_sub_2_io_s_delay_7;
  reg        [376:0]  adder_0_sub_2_io_s_delay_8;
  reg        [376:0]  adder_0_sub_2_io_s_delay_9;
  reg        [376:0]  adder_0_sub_2_io_s_delay_10;
  reg        [376:0]  adder_0_sub_2_io_s_delay_11;
  reg        [376:0]  adder_0_sub_2_io_s_delay_12;
  reg        [376:0]  adder_0_sub_2_io_s_delay_13;
  reg        [376:0]  adder_0_sub_2_io_s_delay_14;
  reg        [376:0]  adder_0_sub_2_io_s_delay_15;
  reg        [376:0]  adder_0_sub_2_io_s_delay_16;
  reg        [376:0]  adder_0_sub_2_io_s_delay_17;
  reg        [376:0]  adder_0_sub_2_io_s_delay_18;
  reg        [376:0]  adder_0_sub_2_io_s_delay_19;
  reg        [376:0]  adder_0_sub_2_io_s_delay_20;
  reg        [376:0]  adder_0_sub_2_io_s_delay_21;
  reg        [376:0]  adder_0_sub_2_io_s_delay_22;
  reg        [376:0]  adder_0_sub_2_io_s_delay_23;
  reg        [376:0]  adder_0_sub_2_io_s_delay_24;
  reg        [376:0]  adder_0_sub_2_io_s_delay_25;
  reg        [376:0]  adder_0_sub_2_io_s_delay_26;
  reg        [376:0]  adder_0_sub_2_io_s_delay_27;
  reg        [376:0]  adder_0_sub_2_io_s_delay_28;
  reg        [376:0]  adder_0_sub_2_io_s_delay_29;
  reg        [376:0]  adder_0_sub_2_io_s_delay_30;
  reg        [376:0]  adder_0_sub_2_io_s_delay_31;
  reg        [376:0]  adder_0_sub_2_io_s_delay_32;
  reg        [376:0]  adder_0_sub_2_io_s_delay_33;
  reg        [376:0]  adder_0_sub_2_io_s_delay_34;
  reg        [376:0]  adder_0_sub_2_io_s_delay_35;
  reg        [376:0]  adder_0_sub_2_io_s_delay_36;
  reg        [376:0]  adder_0_sub_2_io_s_delay_37;
  reg        [376:0]  adder_0_sub_2_io_s_delay_38;
  reg        [376:0]  adder_0_sub_2_io_s_delay_39;
  reg        [376:0]  adder_0_sub_2_io_s_delay_40;
  reg        [376:0]  adder_0_sub_2_io_s_delay_41;
  reg        [376:0]  adder_0_sub_2_io_s_delay_42;
  reg        [376:0]  adder_0_sub_2_io_s_delay_43;
  reg        [376:0]  adder_0_sub_2_io_s_delay_44;
  reg        [376:0]  adder_0_sub_2_io_s_delay_45;
  reg        [376:0]  adder_0_sub_2_io_s_delay_46;
  reg        [376:0]  adder_0_sub_2_io_s_delay_47;
  reg        [376:0]  adder_0_sub_2_io_s_delay_48;
  reg        [376:0]  adder_0_sub_2_io_s_delay_49;
  reg        [376:0]  adder_0_sub_2_io_s_delay_50;
  reg        [376:0]  adder_0_sub_2_io_s_delay_51;
  reg        [376:0]  adder_0_sub_2_io_s_delay_52;
  reg        [376:0]  adder_0_sub_2_io_s_delay_53;
  reg        [376:0]  adder_0_sub_2_io_s_delay_54;
  reg        [376:0]  adder_0_sub_2_io_s_delay_55;
  reg        [376:0]  adder_0_sub_2_io_s_delay_56;
  reg        [376:0]  adder_0_sub_2_io_s_delay_57;
  reg        [376:0]  adder_0_sub_2_io_s_delay_58;
  reg        [376:0]  adder_0_sub_2_io_s_delay_59;
  reg        [376:0]  adder_0_sub_2_io_s_delay_60;
  reg        [376:0]  adder_0_sub_2_io_s_delay_61;
  reg        [376:0]  adder_0_sub_2_io_s_delay_62;
  reg        [376:0]  adder_0_sub_2_io_s_delay_63;
  reg        [376:0]  adder_0_sub_2_io_s_delay_64;
  reg        [376:0]  adder_0_sub_2_io_s_delay_65;
  reg        [376:0]  adder_0_sub_2_io_s_delay_66;
  reg        [376:0]  adder_0_sub_2_io_s_delay_67;
  reg        [376:0]  adder_0_sub_2_io_s_delay_68;
  reg        [376:0]  adder_0_sub_2_io_s_delay_69;
  reg        [376:0]  adder_0_sub_2_io_s_delay_70;
  reg        [376:0]  adder_0_sub_2_io_s_delay_71;
  reg        [376:0]  adder_0_sub_2_io_s_delay_72;
  reg        [376:0]  adder_0_sub_2_io_s_delay_73;
  reg        [376:0]  adder_0_sub_2_io_s_delay_74;
  reg        [376:0]  adder_0_sub_2_io_s_delay_75;
  reg        [376:0]  R9;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_1;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_2;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_3;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_4;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_5;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_6;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_7;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_8;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_9;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_10;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_11;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_12;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_13;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_14;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_15;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_16;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_17;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_18;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_19;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_20;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_21;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_22;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_23;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_24;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_25;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_26;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_27;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_28;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_29;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_30;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_31;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_32;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_33;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_34;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_35;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_36;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_37;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_38;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_39;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_40;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_41;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_42;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_43;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_44;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_45;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_46;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_47;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_48;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_49;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_50;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_51;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_52;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_53;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_54;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_55;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_56;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_57;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_58;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_59;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_60;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_61;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_62;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_63;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_64;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_65;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_66;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_67;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_68;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_69;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_70;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_71;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_72;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_73;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_74;
  reg        [376:0]  adder_0_add_3_1_io_s_delay_75;
  reg        [376:0]  R12;

  KaratsubaMMUL_9 mul_0 (
    .io_a   (sub_0_io_s[376:0]), //i
    .io_b   (sub_1_io_s[376:0]), //i
    .io_p   (mul_0_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL_9 mul_1 (
    .io_a   (add_0_io_s[376:0]  ), //i
    .io_b   (add_1_1_io_s[376:0]), //i
    .io_p   (mul_1_io_p[376:0]  ), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  KaratsubaMMUL_9 mul_2 (
    .io_a   (io_a_T_delay_84[376:0]), //i
    .io_b   (cMul_io_p[376:0]      ), //i
    .io_p   (mul_2_io_p[376:0]     ), //o
    .clk    (clk                   ), //i
    .resetn (resetn                )  //i
  );
  KaratsubaMMUL_9 mul_3 (
    .io_a   (io_a_Z[376:0]    ), //i
    .io_b   (io_b_Z[376:0]    ), //i
    .io_p   (mul_3_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL_9 mul_4 (
    .io_a   (R9[376:0]        ), //i
    .io_b   (sub_3_io_s[376:0]), //i
    .io_p   (mul_4_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL_9 mul_5 (
    .io_a   (add_2_1_io_s[376:0]), //i
    .io_b   (R12[376:0]         ), //i
    .io_p   (mul_5_io_p[376:0]  ), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  KaratsubaMMUL_9 mul_6 (
    .io_a   (sub_3_io_s[376:0]  ), //i
    .io_b   (add_2_1_io_s[376:0]), //i
    .io_p   (mul_6_io_p[376:0]  ), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  KaratsubaMMUL_9 mul_7 (
    .io_a   (R9[376:0]        ), //i
    .io_b   (R12[376:0]       ), //i
    .io_p   (mul_7_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL_9 cMul (
    .io_a   (io_b_T[376:0]                                                                                       ), //i
    .io_b   (377'h196bab03169a4f2ca0b7670ae65fc7437786998c1a32d217f165b2fe0b32139735d947870e3d3e4e02c125684d6e016), //i
    .io_p   (cMul_io_p[376:0]                                                                                    ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  MADD_8 add_0 (
    .io_a   (io_a_Y[376:0]    ), //i
    .io_b   (io_a_X[376:0]    ), //i
    .io_s   (add_0_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_8 add_1_1 (
    .io_a   (io_b_Y[376:0]      ), //i
    .io_b   (io_b_X[376:0]      ), //i
    .io_s   (add_1_1_io_s[376:0]), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  MADD_8 add_2_1 (
    .io_a   (R8[376:0]          ), //i
    .io_b   (mul_2_io_p[376:0]  ), //i
    .io_s   (add_2_1_io_s[376:0]), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  MADD_8 add_3_1 (
    .io_a   (mul_1_io_p[376:0]  ), //i
    .io_b   (mul_0_io_p[376:0]  ), //i
    .io_s   (add_3_1_io_s[376:0]), //o
    .clk    (clk                ), //i
    .resetn (resetn             )  //i
  );
  MADD_12 sub_0 (
    .io_a   (io_a_Y[376:0]    ), //i
    .io_b   (io_a_X[376:0]    ), //i
    .io_s   (sub_0_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_12 sub_1 (
    .io_a   (io_b_Y[376:0]    ), //i
    .io_b   (io_b_X[376:0]    ), //i
    .io_s   (sub_1_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_12 sub_2 (
    .io_a   (mul_1_io_p[376:0]), //i
    .io_b   (mul_0_io_p[376:0]), //i
    .io_s   (sub_2_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_12 sub_3 (
    .io_a   (R8[376:0]        ), //i
    .io_b   (mul_2_io_p[376:0]), //i
    .io_s   (sub_3_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  FineReduction_1 reduction (
    .io_a   (reduction_io_a[377:0]), //i
    .io_r   (reduction_io_r[376:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign reduction_io_a = ({1'd0,mul_3_io_p} <<< 1);
  assign io_s_X = mul_4_io_p;
  assign io_s_Y = mul_5_io_p;
  assign io_s_Z = mul_6_io_p;
  assign io_s_T = mul_7_io_p;
  always @(posedge clk) begin
    io_a_T_delay_1 <= io_a_T;
    io_a_T_delay_2 <= io_a_T_delay_1;
    io_a_T_delay_3 <= io_a_T_delay_2;
    io_a_T_delay_4 <= io_a_T_delay_3;
    io_a_T_delay_5 <= io_a_T_delay_4;
    io_a_T_delay_6 <= io_a_T_delay_5;
    io_a_T_delay_7 <= io_a_T_delay_6;
    io_a_T_delay_8 <= io_a_T_delay_7;
    io_a_T_delay_9 <= io_a_T_delay_8;
    io_a_T_delay_10 <= io_a_T_delay_9;
    io_a_T_delay_11 <= io_a_T_delay_10;
    io_a_T_delay_12 <= io_a_T_delay_11;
    io_a_T_delay_13 <= io_a_T_delay_12;
    io_a_T_delay_14 <= io_a_T_delay_13;
    io_a_T_delay_15 <= io_a_T_delay_14;
    io_a_T_delay_16 <= io_a_T_delay_15;
    io_a_T_delay_17 <= io_a_T_delay_16;
    io_a_T_delay_18 <= io_a_T_delay_17;
    io_a_T_delay_19 <= io_a_T_delay_18;
    io_a_T_delay_20 <= io_a_T_delay_19;
    io_a_T_delay_21 <= io_a_T_delay_20;
    io_a_T_delay_22 <= io_a_T_delay_21;
    io_a_T_delay_23 <= io_a_T_delay_22;
    io_a_T_delay_24 <= io_a_T_delay_23;
    io_a_T_delay_25 <= io_a_T_delay_24;
    io_a_T_delay_26 <= io_a_T_delay_25;
    io_a_T_delay_27 <= io_a_T_delay_26;
    io_a_T_delay_28 <= io_a_T_delay_27;
    io_a_T_delay_29 <= io_a_T_delay_28;
    io_a_T_delay_30 <= io_a_T_delay_29;
    io_a_T_delay_31 <= io_a_T_delay_30;
    io_a_T_delay_32 <= io_a_T_delay_31;
    io_a_T_delay_33 <= io_a_T_delay_32;
    io_a_T_delay_34 <= io_a_T_delay_33;
    io_a_T_delay_35 <= io_a_T_delay_34;
    io_a_T_delay_36 <= io_a_T_delay_35;
    io_a_T_delay_37 <= io_a_T_delay_36;
    io_a_T_delay_38 <= io_a_T_delay_37;
    io_a_T_delay_39 <= io_a_T_delay_38;
    io_a_T_delay_40 <= io_a_T_delay_39;
    io_a_T_delay_41 <= io_a_T_delay_40;
    io_a_T_delay_42 <= io_a_T_delay_41;
    io_a_T_delay_43 <= io_a_T_delay_42;
    io_a_T_delay_44 <= io_a_T_delay_43;
    io_a_T_delay_45 <= io_a_T_delay_44;
    io_a_T_delay_46 <= io_a_T_delay_45;
    io_a_T_delay_47 <= io_a_T_delay_46;
    io_a_T_delay_48 <= io_a_T_delay_47;
    io_a_T_delay_49 <= io_a_T_delay_48;
    io_a_T_delay_50 <= io_a_T_delay_49;
    io_a_T_delay_51 <= io_a_T_delay_50;
    io_a_T_delay_52 <= io_a_T_delay_51;
    io_a_T_delay_53 <= io_a_T_delay_52;
    io_a_T_delay_54 <= io_a_T_delay_53;
    io_a_T_delay_55 <= io_a_T_delay_54;
    io_a_T_delay_56 <= io_a_T_delay_55;
    io_a_T_delay_57 <= io_a_T_delay_56;
    io_a_T_delay_58 <= io_a_T_delay_57;
    io_a_T_delay_59 <= io_a_T_delay_58;
    io_a_T_delay_60 <= io_a_T_delay_59;
    io_a_T_delay_61 <= io_a_T_delay_60;
    io_a_T_delay_62 <= io_a_T_delay_61;
    io_a_T_delay_63 <= io_a_T_delay_62;
    io_a_T_delay_64 <= io_a_T_delay_63;
    io_a_T_delay_65 <= io_a_T_delay_64;
    io_a_T_delay_66 <= io_a_T_delay_65;
    io_a_T_delay_67 <= io_a_T_delay_66;
    io_a_T_delay_68 <= io_a_T_delay_67;
    io_a_T_delay_69 <= io_a_T_delay_68;
    io_a_T_delay_70 <= io_a_T_delay_69;
    io_a_T_delay_71 <= io_a_T_delay_70;
    io_a_T_delay_72 <= io_a_T_delay_71;
    io_a_T_delay_73 <= io_a_T_delay_72;
    io_a_T_delay_74 <= io_a_T_delay_73;
    io_a_T_delay_75 <= io_a_T_delay_74;
    io_a_T_delay_76 <= io_a_T_delay_75;
    io_a_T_delay_77 <= io_a_T_delay_76;
    io_a_T_delay_78 <= io_a_T_delay_77;
    io_a_T_delay_79 <= io_a_T_delay_78;
    io_a_T_delay_80 <= io_a_T_delay_79;
    io_a_T_delay_81 <= io_a_T_delay_80;
    io_a_T_delay_82 <= io_a_T_delay_81;
    io_a_T_delay_83 <= io_a_T_delay_82;
    io_a_T_delay_84 <= io_a_T_delay_83;
    adder_0_reduction_io_r_delay_1 <= reduction_io_r;
    adder_0_reduction_io_r_delay_2 <= adder_0_reduction_io_r_delay_1;
    adder_0_reduction_io_r_delay_3 <= adder_0_reduction_io_r_delay_2;
    adder_0_reduction_io_r_delay_4 <= adder_0_reduction_io_r_delay_3;
    adder_0_reduction_io_r_delay_5 <= adder_0_reduction_io_r_delay_4;
    adder_0_reduction_io_r_delay_6 <= adder_0_reduction_io_r_delay_5;
    adder_0_reduction_io_r_delay_7 <= adder_0_reduction_io_r_delay_6;
    adder_0_reduction_io_r_delay_8 <= adder_0_reduction_io_r_delay_7;
    adder_0_reduction_io_r_delay_9 <= adder_0_reduction_io_r_delay_8;
    adder_0_reduction_io_r_delay_10 <= adder_0_reduction_io_r_delay_9;
    adder_0_reduction_io_r_delay_11 <= adder_0_reduction_io_r_delay_10;
    adder_0_reduction_io_r_delay_12 <= adder_0_reduction_io_r_delay_11;
    adder_0_reduction_io_r_delay_13 <= adder_0_reduction_io_r_delay_12;
    adder_0_reduction_io_r_delay_14 <= adder_0_reduction_io_r_delay_13;
    adder_0_reduction_io_r_delay_15 <= adder_0_reduction_io_r_delay_14;
    adder_0_reduction_io_r_delay_16 <= adder_0_reduction_io_r_delay_15;
    adder_0_reduction_io_r_delay_17 <= adder_0_reduction_io_r_delay_16;
    adder_0_reduction_io_r_delay_18 <= adder_0_reduction_io_r_delay_17;
    adder_0_reduction_io_r_delay_19 <= adder_0_reduction_io_r_delay_18;
    adder_0_reduction_io_r_delay_20 <= adder_0_reduction_io_r_delay_19;
    adder_0_reduction_io_r_delay_21 <= adder_0_reduction_io_r_delay_20;
    adder_0_reduction_io_r_delay_22 <= adder_0_reduction_io_r_delay_21;
    adder_0_reduction_io_r_delay_23 <= adder_0_reduction_io_r_delay_22;
    adder_0_reduction_io_r_delay_24 <= adder_0_reduction_io_r_delay_23;
    adder_0_reduction_io_r_delay_25 <= adder_0_reduction_io_r_delay_24;
    adder_0_reduction_io_r_delay_26 <= adder_0_reduction_io_r_delay_25;
    adder_0_reduction_io_r_delay_27 <= adder_0_reduction_io_r_delay_26;
    adder_0_reduction_io_r_delay_28 <= adder_0_reduction_io_r_delay_27;
    adder_0_reduction_io_r_delay_29 <= adder_0_reduction_io_r_delay_28;
    adder_0_reduction_io_r_delay_30 <= adder_0_reduction_io_r_delay_29;
    adder_0_reduction_io_r_delay_31 <= adder_0_reduction_io_r_delay_30;
    adder_0_reduction_io_r_delay_32 <= adder_0_reduction_io_r_delay_31;
    adder_0_reduction_io_r_delay_33 <= adder_0_reduction_io_r_delay_32;
    adder_0_reduction_io_r_delay_34 <= adder_0_reduction_io_r_delay_33;
    adder_0_reduction_io_r_delay_35 <= adder_0_reduction_io_r_delay_34;
    adder_0_reduction_io_r_delay_36 <= adder_0_reduction_io_r_delay_35;
    adder_0_reduction_io_r_delay_37 <= adder_0_reduction_io_r_delay_36;
    adder_0_reduction_io_r_delay_38 <= adder_0_reduction_io_r_delay_37;
    adder_0_reduction_io_r_delay_39 <= adder_0_reduction_io_r_delay_38;
    adder_0_reduction_io_r_delay_40 <= adder_0_reduction_io_r_delay_39;
    adder_0_reduction_io_r_delay_41 <= adder_0_reduction_io_r_delay_40;
    adder_0_reduction_io_r_delay_42 <= adder_0_reduction_io_r_delay_41;
    adder_0_reduction_io_r_delay_43 <= adder_0_reduction_io_r_delay_42;
    adder_0_reduction_io_r_delay_44 <= adder_0_reduction_io_r_delay_43;
    adder_0_reduction_io_r_delay_45 <= adder_0_reduction_io_r_delay_44;
    adder_0_reduction_io_r_delay_46 <= adder_0_reduction_io_r_delay_45;
    adder_0_reduction_io_r_delay_47 <= adder_0_reduction_io_r_delay_46;
    adder_0_reduction_io_r_delay_48 <= adder_0_reduction_io_r_delay_47;
    adder_0_reduction_io_r_delay_49 <= adder_0_reduction_io_r_delay_48;
    adder_0_reduction_io_r_delay_50 <= adder_0_reduction_io_r_delay_49;
    adder_0_reduction_io_r_delay_51 <= adder_0_reduction_io_r_delay_50;
    adder_0_reduction_io_r_delay_52 <= adder_0_reduction_io_r_delay_51;
    adder_0_reduction_io_r_delay_53 <= adder_0_reduction_io_r_delay_52;
    adder_0_reduction_io_r_delay_54 <= adder_0_reduction_io_r_delay_53;
    adder_0_reduction_io_r_delay_55 <= adder_0_reduction_io_r_delay_54;
    adder_0_reduction_io_r_delay_56 <= adder_0_reduction_io_r_delay_55;
    adder_0_reduction_io_r_delay_57 <= adder_0_reduction_io_r_delay_56;
    adder_0_reduction_io_r_delay_58 <= adder_0_reduction_io_r_delay_57;
    adder_0_reduction_io_r_delay_59 <= adder_0_reduction_io_r_delay_58;
    adder_0_reduction_io_r_delay_60 <= adder_0_reduction_io_r_delay_59;
    adder_0_reduction_io_r_delay_61 <= adder_0_reduction_io_r_delay_60;
    adder_0_reduction_io_r_delay_62 <= adder_0_reduction_io_r_delay_61;
    adder_0_reduction_io_r_delay_63 <= adder_0_reduction_io_r_delay_62;
    adder_0_reduction_io_r_delay_64 <= adder_0_reduction_io_r_delay_63;
    adder_0_reduction_io_r_delay_65 <= adder_0_reduction_io_r_delay_64;
    adder_0_reduction_io_r_delay_66 <= adder_0_reduction_io_r_delay_65;
    adder_0_reduction_io_r_delay_67 <= adder_0_reduction_io_r_delay_66;
    adder_0_reduction_io_r_delay_68 <= adder_0_reduction_io_r_delay_67;
    adder_0_reduction_io_r_delay_69 <= adder_0_reduction_io_r_delay_68;
    adder_0_reduction_io_r_delay_70 <= adder_0_reduction_io_r_delay_69;
    adder_0_reduction_io_r_delay_71 <= adder_0_reduction_io_r_delay_70;
    adder_0_reduction_io_r_delay_72 <= adder_0_reduction_io_r_delay_71;
    adder_0_reduction_io_r_delay_73 <= adder_0_reduction_io_r_delay_72;
    adder_0_reduction_io_r_delay_74 <= adder_0_reduction_io_r_delay_73;
    adder_0_reduction_io_r_delay_75 <= adder_0_reduction_io_r_delay_74;
    adder_0_reduction_io_r_delay_76 <= adder_0_reduction_io_r_delay_75;
    R8 <= adder_0_reduction_io_r_delay_76;
    adder_0_sub_2_io_s_delay_1 <= sub_2_io_s;
    adder_0_sub_2_io_s_delay_2 <= adder_0_sub_2_io_s_delay_1;
    adder_0_sub_2_io_s_delay_3 <= adder_0_sub_2_io_s_delay_2;
    adder_0_sub_2_io_s_delay_4 <= adder_0_sub_2_io_s_delay_3;
    adder_0_sub_2_io_s_delay_5 <= adder_0_sub_2_io_s_delay_4;
    adder_0_sub_2_io_s_delay_6 <= adder_0_sub_2_io_s_delay_5;
    adder_0_sub_2_io_s_delay_7 <= adder_0_sub_2_io_s_delay_6;
    adder_0_sub_2_io_s_delay_8 <= adder_0_sub_2_io_s_delay_7;
    adder_0_sub_2_io_s_delay_9 <= adder_0_sub_2_io_s_delay_8;
    adder_0_sub_2_io_s_delay_10 <= adder_0_sub_2_io_s_delay_9;
    adder_0_sub_2_io_s_delay_11 <= adder_0_sub_2_io_s_delay_10;
    adder_0_sub_2_io_s_delay_12 <= adder_0_sub_2_io_s_delay_11;
    adder_0_sub_2_io_s_delay_13 <= adder_0_sub_2_io_s_delay_12;
    adder_0_sub_2_io_s_delay_14 <= adder_0_sub_2_io_s_delay_13;
    adder_0_sub_2_io_s_delay_15 <= adder_0_sub_2_io_s_delay_14;
    adder_0_sub_2_io_s_delay_16 <= adder_0_sub_2_io_s_delay_15;
    adder_0_sub_2_io_s_delay_17 <= adder_0_sub_2_io_s_delay_16;
    adder_0_sub_2_io_s_delay_18 <= adder_0_sub_2_io_s_delay_17;
    adder_0_sub_2_io_s_delay_19 <= adder_0_sub_2_io_s_delay_18;
    adder_0_sub_2_io_s_delay_20 <= adder_0_sub_2_io_s_delay_19;
    adder_0_sub_2_io_s_delay_21 <= adder_0_sub_2_io_s_delay_20;
    adder_0_sub_2_io_s_delay_22 <= adder_0_sub_2_io_s_delay_21;
    adder_0_sub_2_io_s_delay_23 <= adder_0_sub_2_io_s_delay_22;
    adder_0_sub_2_io_s_delay_24 <= adder_0_sub_2_io_s_delay_23;
    adder_0_sub_2_io_s_delay_25 <= adder_0_sub_2_io_s_delay_24;
    adder_0_sub_2_io_s_delay_26 <= adder_0_sub_2_io_s_delay_25;
    adder_0_sub_2_io_s_delay_27 <= adder_0_sub_2_io_s_delay_26;
    adder_0_sub_2_io_s_delay_28 <= adder_0_sub_2_io_s_delay_27;
    adder_0_sub_2_io_s_delay_29 <= adder_0_sub_2_io_s_delay_28;
    adder_0_sub_2_io_s_delay_30 <= adder_0_sub_2_io_s_delay_29;
    adder_0_sub_2_io_s_delay_31 <= adder_0_sub_2_io_s_delay_30;
    adder_0_sub_2_io_s_delay_32 <= adder_0_sub_2_io_s_delay_31;
    adder_0_sub_2_io_s_delay_33 <= adder_0_sub_2_io_s_delay_32;
    adder_0_sub_2_io_s_delay_34 <= adder_0_sub_2_io_s_delay_33;
    adder_0_sub_2_io_s_delay_35 <= adder_0_sub_2_io_s_delay_34;
    adder_0_sub_2_io_s_delay_36 <= adder_0_sub_2_io_s_delay_35;
    adder_0_sub_2_io_s_delay_37 <= adder_0_sub_2_io_s_delay_36;
    adder_0_sub_2_io_s_delay_38 <= adder_0_sub_2_io_s_delay_37;
    adder_0_sub_2_io_s_delay_39 <= adder_0_sub_2_io_s_delay_38;
    adder_0_sub_2_io_s_delay_40 <= adder_0_sub_2_io_s_delay_39;
    adder_0_sub_2_io_s_delay_41 <= adder_0_sub_2_io_s_delay_40;
    adder_0_sub_2_io_s_delay_42 <= adder_0_sub_2_io_s_delay_41;
    adder_0_sub_2_io_s_delay_43 <= adder_0_sub_2_io_s_delay_42;
    adder_0_sub_2_io_s_delay_44 <= adder_0_sub_2_io_s_delay_43;
    adder_0_sub_2_io_s_delay_45 <= adder_0_sub_2_io_s_delay_44;
    adder_0_sub_2_io_s_delay_46 <= adder_0_sub_2_io_s_delay_45;
    adder_0_sub_2_io_s_delay_47 <= adder_0_sub_2_io_s_delay_46;
    adder_0_sub_2_io_s_delay_48 <= adder_0_sub_2_io_s_delay_47;
    adder_0_sub_2_io_s_delay_49 <= adder_0_sub_2_io_s_delay_48;
    adder_0_sub_2_io_s_delay_50 <= adder_0_sub_2_io_s_delay_49;
    adder_0_sub_2_io_s_delay_51 <= adder_0_sub_2_io_s_delay_50;
    adder_0_sub_2_io_s_delay_52 <= adder_0_sub_2_io_s_delay_51;
    adder_0_sub_2_io_s_delay_53 <= adder_0_sub_2_io_s_delay_52;
    adder_0_sub_2_io_s_delay_54 <= adder_0_sub_2_io_s_delay_53;
    adder_0_sub_2_io_s_delay_55 <= adder_0_sub_2_io_s_delay_54;
    adder_0_sub_2_io_s_delay_56 <= adder_0_sub_2_io_s_delay_55;
    adder_0_sub_2_io_s_delay_57 <= adder_0_sub_2_io_s_delay_56;
    adder_0_sub_2_io_s_delay_58 <= adder_0_sub_2_io_s_delay_57;
    adder_0_sub_2_io_s_delay_59 <= adder_0_sub_2_io_s_delay_58;
    adder_0_sub_2_io_s_delay_60 <= adder_0_sub_2_io_s_delay_59;
    adder_0_sub_2_io_s_delay_61 <= adder_0_sub_2_io_s_delay_60;
    adder_0_sub_2_io_s_delay_62 <= adder_0_sub_2_io_s_delay_61;
    adder_0_sub_2_io_s_delay_63 <= adder_0_sub_2_io_s_delay_62;
    adder_0_sub_2_io_s_delay_64 <= adder_0_sub_2_io_s_delay_63;
    adder_0_sub_2_io_s_delay_65 <= adder_0_sub_2_io_s_delay_64;
    adder_0_sub_2_io_s_delay_66 <= adder_0_sub_2_io_s_delay_65;
    adder_0_sub_2_io_s_delay_67 <= adder_0_sub_2_io_s_delay_66;
    adder_0_sub_2_io_s_delay_68 <= adder_0_sub_2_io_s_delay_67;
    adder_0_sub_2_io_s_delay_69 <= adder_0_sub_2_io_s_delay_68;
    adder_0_sub_2_io_s_delay_70 <= adder_0_sub_2_io_s_delay_69;
    adder_0_sub_2_io_s_delay_71 <= adder_0_sub_2_io_s_delay_70;
    adder_0_sub_2_io_s_delay_72 <= adder_0_sub_2_io_s_delay_71;
    adder_0_sub_2_io_s_delay_73 <= adder_0_sub_2_io_s_delay_72;
    adder_0_sub_2_io_s_delay_74 <= adder_0_sub_2_io_s_delay_73;
    adder_0_sub_2_io_s_delay_75 <= adder_0_sub_2_io_s_delay_74;
    R9 <= adder_0_sub_2_io_s_delay_75;
    adder_0_add_3_1_io_s_delay_1 <= add_3_1_io_s;
    adder_0_add_3_1_io_s_delay_2 <= adder_0_add_3_1_io_s_delay_1;
    adder_0_add_3_1_io_s_delay_3 <= adder_0_add_3_1_io_s_delay_2;
    adder_0_add_3_1_io_s_delay_4 <= adder_0_add_3_1_io_s_delay_3;
    adder_0_add_3_1_io_s_delay_5 <= adder_0_add_3_1_io_s_delay_4;
    adder_0_add_3_1_io_s_delay_6 <= adder_0_add_3_1_io_s_delay_5;
    adder_0_add_3_1_io_s_delay_7 <= adder_0_add_3_1_io_s_delay_6;
    adder_0_add_3_1_io_s_delay_8 <= adder_0_add_3_1_io_s_delay_7;
    adder_0_add_3_1_io_s_delay_9 <= adder_0_add_3_1_io_s_delay_8;
    adder_0_add_3_1_io_s_delay_10 <= adder_0_add_3_1_io_s_delay_9;
    adder_0_add_3_1_io_s_delay_11 <= adder_0_add_3_1_io_s_delay_10;
    adder_0_add_3_1_io_s_delay_12 <= adder_0_add_3_1_io_s_delay_11;
    adder_0_add_3_1_io_s_delay_13 <= adder_0_add_3_1_io_s_delay_12;
    adder_0_add_3_1_io_s_delay_14 <= adder_0_add_3_1_io_s_delay_13;
    adder_0_add_3_1_io_s_delay_15 <= adder_0_add_3_1_io_s_delay_14;
    adder_0_add_3_1_io_s_delay_16 <= adder_0_add_3_1_io_s_delay_15;
    adder_0_add_3_1_io_s_delay_17 <= adder_0_add_3_1_io_s_delay_16;
    adder_0_add_3_1_io_s_delay_18 <= adder_0_add_3_1_io_s_delay_17;
    adder_0_add_3_1_io_s_delay_19 <= adder_0_add_3_1_io_s_delay_18;
    adder_0_add_3_1_io_s_delay_20 <= adder_0_add_3_1_io_s_delay_19;
    adder_0_add_3_1_io_s_delay_21 <= adder_0_add_3_1_io_s_delay_20;
    adder_0_add_3_1_io_s_delay_22 <= adder_0_add_3_1_io_s_delay_21;
    adder_0_add_3_1_io_s_delay_23 <= adder_0_add_3_1_io_s_delay_22;
    adder_0_add_3_1_io_s_delay_24 <= adder_0_add_3_1_io_s_delay_23;
    adder_0_add_3_1_io_s_delay_25 <= adder_0_add_3_1_io_s_delay_24;
    adder_0_add_3_1_io_s_delay_26 <= adder_0_add_3_1_io_s_delay_25;
    adder_0_add_3_1_io_s_delay_27 <= adder_0_add_3_1_io_s_delay_26;
    adder_0_add_3_1_io_s_delay_28 <= adder_0_add_3_1_io_s_delay_27;
    adder_0_add_3_1_io_s_delay_29 <= adder_0_add_3_1_io_s_delay_28;
    adder_0_add_3_1_io_s_delay_30 <= adder_0_add_3_1_io_s_delay_29;
    adder_0_add_3_1_io_s_delay_31 <= adder_0_add_3_1_io_s_delay_30;
    adder_0_add_3_1_io_s_delay_32 <= adder_0_add_3_1_io_s_delay_31;
    adder_0_add_3_1_io_s_delay_33 <= adder_0_add_3_1_io_s_delay_32;
    adder_0_add_3_1_io_s_delay_34 <= adder_0_add_3_1_io_s_delay_33;
    adder_0_add_3_1_io_s_delay_35 <= adder_0_add_3_1_io_s_delay_34;
    adder_0_add_3_1_io_s_delay_36 <= adder_0_add_3_1_io_s_delay_35;
    adder_0_add_3_1_io_s_delay_37 <= adder_0_add_3_1_io_s_delay_36;
    adder_0_add_3_1_io_s_delay_38 <= adder_0_add_3_1_io_s_delay_37;
    adder_0_add_3_1_io_s_delay_39 <= adder_0_add_3_1_io_s_delay_38;
    adder_0_add_3_1_io_s_delay_40 <= adder_0_add_3_1_io_s_delay_39;
    adder_0_add_3_1_io_s_delay_41 <= adder_0_add_3_1_io_s_delay_40;
    adder_0_add_3_1_io_s_delay_42 <= adder_0_add_3_1_io_s_delay_41;
    adder_0_add_3_1_io_s_delay_43 <= adder_0_add_3_1_io_s_delay_42;
    adder_0_add_3_1_io_s_delay_44 <= adder_0_add_3_1_io_s_delay_43;
    adder_0_add_3_1_io_s_delay_45 <= adder_0_add_3_1_io_s_delay_44;
    adder_0_add_3_1_io_s_delay_46 <= adder_0_add_3_1_io_s_delay_45;
    adder_0_add_3_1_io_s_delay_47 <= adder_0_add_3_1_io_s_delay_46;
    adder_0_add_3_1_io_s_delay_48 <= adder_0_add_3_1_io_s_delay_47;
    adder_0_add_3_1_io_s_delay_49 <= adder_0_add_3_1_io_s_delay_48;
    adder_0_add_3_1_io_s_delay_50 <= adder_0_add_3_1_io_s_delay_49;
    adder_0_add_3_1_io_s_delay_51 <= adder_0_add_3_1_io_s_delay_50;
    adder_0_add_3_1_io_s_delay_52 <= adder_0_add_3_1_io_s_delay_51;
    adder_0_add_3_1_io_s_delay_53 <= adder_0_add_3_1_io_s_delay_52;
    adder_0_add_3_1_io_s_delay_54 <= adder_0_add_3_1_io_s_delay_53;
    adder_0_add_3_1_io_s_delay_55 <= adder_0_add_3_1_io_s_delay_54;
    adder_0_add_3_1_io_s_delay_56 <= adder_0_add_3_1_io_s_delay_55;
    adder_0_add_3_1_io_s_delay_57 <= adder_0_add_3_1_io_s_delay_56;
    adder_0_add_3_1_io_s_delay_58 <= adder_0_add_3_1_io_s_delay_57;
    adder_0_add_3_1_io_s_delay_59 <= adder_0_add_3_1_io_s_delay_58;
    adder_0_add_3_1_io_s_delay_60 <= adder_0_add_3_1_io_s_delay_59;
    adder_0_add_3_1_io_s_delay_61 <= adder_0_add_3_1_io_s_delay_60;
    adder_0_add_3_1_io_s_delay_62 <= adder_0_add_3_1_io_s_delay_61;
    adder_0_add_3_1_io_s_delay_63 <= adder_0_add_3_1_io_s_delay_62;
    adder_0_add_3_1_io_s_delay_64 <= adder_0_add_3_1_io_s_delay_63;
    adder_0_add_3_1_io_s_delay_65 <= adder_0_add_3_1_io_s_delay_64;
    adder_0_add_3_1_io_s_delay_66 <= adder_0_add_3_1_io_s_delay_65;
    adder_0_add_3_1_io_s_delay_67 <= adder_0_add_3_1_io_s_delay_66;
    adder_0_add_3_1_io_s_delay_68 <= adder_0_add_3_1_io_s_delay_67;
    adder_0_add_3_1_io_s_delay_69 <= adder_0_add_3_1_io_s_delay_68;
    adder_0_add_3_1_io_s_delay_70 <= adder_0_add_3_1_io_s_delay_69;
    adder_0_add_3_1_io_s_delay_71 <= adder_0_add_3_1_io_s_delay_70;
    adder_0_add_3_1_io_s_delay_72 <= adder_0_add_3_1_io_s_delay_71;
    adder_0_add_3_1_io_s_delay_73 <= adder_0_add_3_1_io_s_delay_72;
    adder_0_add_3_1_io_s_delay_74 <= adder_0_add_3_1_io_s_delay_73;
    adder_0_add_3_1_io_s_delay_75 <= adder_0_add_3_1_io_s_delay_74;
    R12 <= adder_0_add_3_1_io_s_delay_75;
  end


endmodule

//DWSRFIFO_1 replaced by DWSRFIFO

module DWSRFIFO (
  input               io_dataIn_0_valid,
  input      [376:0]  io_dataIn_0_payload_a_X,
  input      [376:0]  io_dataIn_0_payload_a_Y,
  input      [376:0]  io_dataIn_0_payload_a_Z,
  input      [376:0]  io_dataIn_0_payload_a_T,
  input      [376:0]  io_dataIn_0_payload_b_X,
  input      [376:0]  io_dataIn_0_payload_b_Y,
  input      [376:0]  io_dataIn_0_payload_b_Z,
  input      [376:0]  io_dataIn_0_payload_b_T,
  input      [15:0]   io_dataIn_0_payload_address,
  input               io_dataIn_1_valid,
  input      [376:0]  io_dataIn_1_payload_a_X,
  input      [376:0]  io_dataIn_1_payload_a_Y,
  input      [376:0]  io_dataIn_1_payload_a_Z,
  input      [376:0]  io_dataIn_1_payload_a_T,
  input      [376:0]  io_dataIn_1_payload_b_X,
  input      [376:0]  io_dataIn_1_payload_b_Y,
  input      [376:0]  io_dataIn_1_payload_b_Z,
  input      [376:0]  io_dataIn_1_payload_b_T,
  input      [15:0]   io_dataIn_1_payload_address,
  output              io_dataOut_valid,
  output     [376:0]  io_dataOut_payload_a_X,
  output     [376:0]  io_dataOut_payload_a_Y,
  output     [376:0]  io_dataOut_payload_a_Z,
  output     [376:0]  io_dataOut_payload_a_T,
  output     [376:0]  io_dataOut_payload_b_X,
  output     [376:0]  io_dataOut_payload_b_Y,
  output     [376:0]  io_dataOut_payload_b_Z,
  output     [376:0]  io_dataOut_payload_b_T,
  output     [15:0]   io_dataOut_payload_address,
  input               clk,
  input               resetn
);

  wire       [376:0]  ram_io_rData_a_X;
  wire       [376:0]  ram_io_rData_a_Y;
  wire       [376:0]  ram_io_rData_a_Z;
  wire       [376:0]  ram_io_rData_a_T;
  wire       [376:0]  ram_io_rData_b_X;
  wire       [376:0]  ram_io_rData_b_Y;
  wire       [376:0]  ram_io_rData_b_Z;
  wire       [376:0]  ram_io_rData_b_T;
  wire       [15:0]   ram_io_rData_address;
  wire       [7:0]    _zz_pushPtr_valueNext;
  wire       [0:0]    _zz_pushPtr_valueNext_1;
  wire       [7:0]    _zz_popPtr_valueNext;
  wire       [0:0]    _zz_popPtr_valueNext_1;
  reg                 pushPtr_willIncrement;
  wire                pushPtr_willClear;
  reg        [7:0]    pushPtr_valueNext;
  reg        [7:0]    pushPtr_value;
  reg                 pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  wire                popPtr_willClear;
  reg        [7:0]    popPtr_valueNext;
  reg        [7:0]    popPtr_value;
  reg                 popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  reg                 empty;
  reg                 _zz_io_dataOut_valid;
  reg                 _zz_io_dataOut_valid_1;
  reg                 _zz_io_dataOut_valid_2;
  reg                 _zz_io_dataOut_valid_3;
  reg                 io_dataIn_1_valid_delay_1;
  reg                 io_dataIn_1_valid_delay_2;
  reg                 io_dataIn_1_valid_delay_3;
  reg                 io_dataIn_1_valid_delay_4;
  reg        [376:0]  io_dataIn_1_payload_delay_1_a_X;
  reg        [376:0]  io_dataIn_1_payload_delay_1_a_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_1_a_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_1_a_T;
  reg        [376:0]  io_dataIn_1_payload_delay_1_b_X;
  reg        [376:0]  io_dataIn_1_payload_delay_1_b_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_1_b_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_1_b_T;
  reg        [15:0]   io_dataIn_1_payload_delay_1_address;
  reg        [376:0]  io_dataIn_1_payload_delay_2_a_X;
  reg        [376:0]  io_dataIn_1_payload_delay_2_a_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_2_a_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_2_a_T;
  reg        [376:0]  io_dataIn_1_payload_delay_2_b_X;
  reg        [376:0]  io_dataIn_1_payload_delay_2_b_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_2_b_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_2_b_T;
  reg        [15:0]   io_dataIn_1_payload_delay_2_address;
  reg        [376:0]  io_dataIn_1_payload_delay_3_a_X;
  reg        [376:0]  io_dataIn_1_payload_delay_3_a_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_3_a_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_3_a_T;
  reg        [376:0]  io_dataIn_1_payload_delay_3_b_X;
  reg        [376:0]  io_dataIn_1_payload_delay_3_b_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_3_b_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_3_b_T;
  reg        [15:0]   io_dataIn_1_payload_delay_3_address;
  reg        [376:0]  io_dataIn_1_payload_delay_4_a_X;
  reg        [376:0]  io_dataIn_1_payload_delay_4_a_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_4_a_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_4_a_T;
  reg        [376:0]  io_dataIn_1_payload_delay_4_b_X;
  reg        [376:0]  io_dataIn_1_payload_delay_4_b_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_4_b_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_4_b_T;
  reg        [15:0]   io_dataIn_1_payload_delay_4_address;
  wire                when_DWSRFIFO_l41;

  assign _zz_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign _zz_pushPtr_valueNext = {7'd0, _zz_pushPtr_valueNext_1};
  assign _zz_popPtr_valueNext_1 = popPtr_willIncrement;
  assign _zz_popPtr_valueNext = {7'd0, _zz_popPtr_valueNext_1};
  SDPRAM_1 ram (
    .io_we            (io_dataIn_0_valid                ), //i
    .io_wAddress      (pushPtr_value[7:0]               ), //i
    .io_wData_a_X     (io_dataIn_0_payload_a_X[376:0]   ), //i
    .io_wData_a_Y     (io_dataIn_0_payload_a_Y[376:0]   ), //i
    .io_wData_a_Z     (io_dataIn_0_payload_a_Z[376:0]   ), //i
    .io_wData_a_T     (io_dataIn_0_payload_a_T[376:0]   ), //i
    .io_wData_b_X     (io_dataIn_0_payload_b_X[376:0]   ), //i
    .io_wData_b_Y     (io_dataIn_0_payload_b_Y[376:0]   ), //i
    .io_wData_b_Z     (io_dataIn_0_payload_b_Z[376:0]   ), //i
    .io_wData_b_T     (io_dataIn_0_payload_b_T[376:0]   ), //i
    .io_wData_address (io_dataIn_0_payload_address[15:0]), //i
    .io_re            (1'b1                             ), //i
    .io_rAddress      (popPtr_value[7:0]                ), //i
    .io_rData_a_X     (ram_io_rData_a_X[376:0]          ), //o
    .io_rData_a_Y     (ram_io_rData_a_Y[376:0]          ), //o
    .io_rData_a_Z     (ram_io_rData_a_Z[376:0]          ), //o
    .io_rData_a_T     (ram_io_rData_a_T[376:0]          ), //o
    .io_rData_b_X     (ram_io_rData_b_X[376:0]          ), //o
    .io_rData_b_Y     (ram_io_rData_b_Y[376:0]          ), //o
    .io_rData_b_Z     (ram_io_rData_b_Z[376:0]          ), //o
    .io_rData_b_T     (ram_io_rData_b_T[376:0]          ), //o
    .io_rData_address (ram_io_rData_address[15:0]       ), //o
    .clk              (clk                              ), //i
    .resetn           (resetn                           )  //i
  );
  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(io_dataIn_0_valid) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  assign pushPtr_willClear = 1'b0;
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    pushPtr_valueNext = (pushPtr_value + _zz_pushPtr_valueNext);
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 8'h0;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(when_DWSRFIFO_l41) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  assign popPtr_willClear = 1'b0;
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    popPtr_valueNext = (popPtr_value + _zz_popPtr_valueNext);
    if(popPtr_willClear) begin
      popPtr_valueNext = 8'h0;
    end
  end

  assign io_dataOut_valid = _zz_io_dataOut_valid_3;
  assign io_dataOut_payload_a_X = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_a_X : ram_io_rData_a_X);
  assign io_dataOut_payload_a_Y = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_a_Y : ram_io_rData_a_Y);
  assign io_dataOut_payload_a_Z = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_a_Z : ram_io_rData_a_Z);
  assign io_dataOut_payload_a_T = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_a_T : ram_io_rData_a_T);
  assign io_dataOut_payload_b_X = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_b_X : ram_io_rData_b_X);
  assign io_dataOut_payload_b_Y = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_b_Y : ram_io_rData_b_Y);
  assign io_dataOut_payload_b_Z = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_b_Z : ram_io_rData_b_Z);
  assign io_dataOut_payload_b_T = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_b_T : ram_io_rData_b_T);
  assign io_dataOut_payload_address = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_address : ram_io_rData_address);
  assign when_DWSRFIFO_l41 = ((! empty) && (! io_dataIn_1_valid));
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      pushPtr_value <= 8'h0;
      pushPtr_willOverflowIfInc <= 1'b0;
      popPtr_value <= 8'h0;
      popPtr_willOverflowIfInc <= 1'b0;
      empty <= 1'b1;
      _zz_io_dataOut_valid <= 1'b0;
      _zz_io_dataOut_valid_1 <= 1'b0;
      _zz_io_dataOut_valid_2 <= 1'b0;
      _zz_io_dataOut_valid_3 <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      pushPtr_willOverflowIfInc <= (pushPtr_valueNext == 8'hff);
      popPtr_value <= popPtr_valueNext;
      popPtr_willOverflowIfInc <= (popPtr_valueNext == 8'hff);
      empty <= (pushPtr_value == popPtr_valueNext);
      _zz_io_dataOut_valid <= ((! empty) || io_dataIn_1_valid);
      _zz_io_dataOut_valid_1 <= _zz_io_dataOut_valid;
      _zz_io_dataOut_valid_2 <= _zz_io_dataOut_valid_1;
      _zz_io_dataOut_valid_3 <= _zz_io_dataOut_valid_2;
    end
  end

  always @(posedge clk) begin
    io_dataIn_1_valid_delay_1 <= io_dataIn_1_valid;
    io_dataIn_1_valid_delay_2 <= io_dataIn_1_valid_delay_1;
    io_dataIn_1_valid_delay_3 <= io_dataIn_1_valid_delay_2;
    io_dataIn_1_valid_delay_4 <= io_dataIn_1_valid_delay_3;
    io_dataIn_1_payload_delay_1_a_X <= io_dataIn_1_payload_a_X;
    io_dataIn_1_payload_delay_1_a_Y <= io_dataIn_1_payload_a_Y;
    io_dataIn_1_payload_delay_1_a_Z <= io_dataIn_1_payload_a_Z;
    io_dataIn_1_payload_delay_1_a_T <= io_dataIn_1_payload_a_T;
    io_dataIn_1_payload_delay_1_b_X <= io_dataIn_1_payload_b_X;
    io_dataIn_1_payload_delay_1_b_Y <= io_dataIn_1_payload_b_Y;
    io_dataIn_1_payload_delay_1_b_Z <= io_dataIn_1_payload_b_Z;
    io_dataIn_1_payload_delay_1_b_T <= io_dataIn_1_payload_b_T;
    io_dataIn_1_payload_delay_1_address <= io_dataIn_1_payload_address;
    io_dataIn_1_payload_delay_2_a_X <= io_dataIn_1_payload_delay_1_a_X;
    io_dataIn_1_payload_delay_2_a_Y <= io_dataIn_1_payload_delay_1_a_Y;
    io_dataIn_1_payload_delay_2_a_Z <= io_dataIn_1_payload_delay_1_a_Z;
    io_dataIn_1_payload_delay_2_a_T <= io_dataIn_1_payload_delay_1_a_T;
    io_dataIn_1_payload_delay_2_b_X <= io_dataIn_1_payload_delay_1_b_X;
    io_dataIn_1_payload_delay_2_b_Y <= io_dataIn_1_payload_delay_1_b_Y;
    io_dataIn_1_payload_delay_2_b_Z <= io_dataIn_1_payload_delay_1_b_Z;
    io_dataIn_1_payload_delay_2_b_T <= io_dataIn_1_payload_delay_1_b_T;
    io_dataIn_1_payload_delay_2_address <= io_dataIn_1_payload_delay_1_address;
    io_dataIn_1_payload_delay_3_a_X <= io_dataIn_1_payload_delay_2_a_X;
    io_dataIn_1_payload_delay_3_a_Y <= io_dataIn_1_payload_delay_2_a_Y;
    io_dataIn_1_payload_delay_3_a_Z <= io_dataIn_1_payload_delay_2_a_Z;
    io_dataIn_1_payload_delay_3_a_T <= io_dataIn_1_payload_delay_2_a_T;
    io_dataIn_1_payload_delay_3_b_X <= io_dataIn_1_payload_delay_2_b_X;
    io_dataIn_1_payload_delay_3_b_Y <= io_dataIn_1_payload_delay_2_b_Y;
    io_dataIn_1_payload_delay_3_b_Z <= io_dataIn_1_payload_delay_2_b_Z;
    io_dataIn_1_payload_delay_3_b_T <= io_dataIn_1_payload_delay_2_b_T;
    io_dataIn_1_payload_delay_3_address <= io_dataIn_1_payload_delay_2_address;
    io_dataIn_1_payload_delay_4_a_X <= io_dataIn_1_payload_delay_3_a_X;
    io_dataIn_1_payload_delay_4_a_Y <= io_dataIn_1_payload_delay_3_a_Y;
    io_dataIn_1_payload_delay_4_a_Z <= io_dataIn_1_payload_delay_3_a_Z;
    io_dataIn_1_payload_delay_4_a_T <= io_dataIn_1_payload_delay_3_a_T;
    io_dataIn_1_payload_delay_4_b_X <= io_dataIn_1_payload_delay_3_b_X;
    io_dataIn_1_payload_delay_4_b_Y <= io_dataIn_1_payload_delay_3_b_Y;
    io_dataIn_1_payload_delay_4_b_Z <= io_dataIn_1_payload_delay_3_b_Z;
    io_dataIn_1_payload_delay_4_b_T <= io_dataIn_1_payload_delay_3_b_T;
    io_dataIn_1_payload_delay_4_address <= io_dataIn_1_payload_delay_3_address;
  end


endmodule

//DataRam_1 replaced by DataRam

module DataRam (
  input               io_we_0,
  input               io_we_1,
  input      [15:0]   io_address_0,
  input      [15:0]   io_address_1,
  input      [376:0]  io_wData_0_X,
  input      [376:0]  io_wData_0_Y,
  input      [376:0]  io_wData_0_Z,
  input      [376:0]  io_wData_0_T,
  input      [376:0]  io_wData_1_X,
  input      [376:0]  io_wData_1_Y,
  input      [376:0]  io_wData_1_Z,
  input      [376:0]  io_wData_1_T,
  input               io_state_0,
  input               io_state_1,
  output     [376:0]  io_rData_0_X,
  output     [376:0]  io_rData_0_Y,
  output     [376:0]  io_rData_0_Z,
  output     [376:0]  io_rData_0_T,
  output     [376:0]  io_rData_1_X,
  output     [376:0]  io_rData_1_Y,
  output     [376:0]  io_rData_1_Z,
  output     [376:0]  io_rData_1_T,
  input      [376:0]  io_pInit_X,
  input      [376:0]  io_pInit_Y,
  input      [376:0]  io_pInit_Z,
  input      [376:0]  io_pInit_T,
  input               clk,
  input               resetn
);

  wire       [376:0]  ram_io_rData_0_X;
  wire       [376:0]  ram_io_rData_0_Y;
  wire       [376:0]  ram_io_rData_0_Z;
  wire       [376:0]  ram_io_rData_0_T;
  wire       [376:0]  ram_io_rData_1_X;
  wire       [376:0]  ram_io_rData_1_Y;
  wire       [376:0]  ram_io_rData_1_Z;
  wire       [376:0]  ram_io_rData_1_T;
  reg        [376:0]  _zz_io_rData_0_X;
  reg        [376:0]  _zz_io_rData_0_Y;
  reg        [376:0]  _zz_io_rData_0_Z;
  reg        [376:0]  _zz_io_rData_0_T;
  reg        [376:0]  _zz_io_rData_1_X;
  reg        [376:0]  _zz_io_rData_1_Y;
  reg        [376:0]  _zz_io_rData_1_Z;
  reg        [376:0]  _zz_io_rData_1_T;

  TDPRAM_1 ram (
    .io_we_0      (io_we_0                ), //i
    .io_we_1      (io_we_1                ), //i
    .io_address_0 (io_address_0[15:0]     ), //i
    .io_address_1 (io_address_1[15:0]     ), //i
    .io_wData_0_X (io_wData_0_X[376:0]    ), //i
    .io_wData_0_Y (io_wData_0_Y[376:0]    ), //i
    .io_wData_0_Z (io_wData_0_Z[376:0]    ), //i
    .io_wData_0_T (io_wData_0_T[376:0]    ), //i
    .io_wData_1_X (io_wData_1_X[376:0]    ), //i
    .io_wData_1_Y (io_wData_1_Y[376:0]    ), //i
    .io_wData_1_Z (io_wData_1_Z[376:0]    ), //i
    .io_wData_1_T (io_wData_1_T[376:0]    ), //i
    .io_ce_0      (1'b1                   ), //i
    .io_ce_1      (1'b1                   ), //i
    .io_rData_0_X (ram_io_rData_0_X[376:0]), //o
    .io_rData_0_Y (ram_io_rData_0_Y[376:0]), //o
    .io_rData_0_Z (ram_io_rData_0_Z[376:0]), //o
    .io_rData_0_T (ram_io_rData_0_T[376:0]), //o
    .io_rData_1_X (ram_io_rData_1_X[376:0]), //o
    .io_rData_1_Y (ram_io_rData_1_Y[376:0]), //o
    .io_rData_1_Z (ram_io_rData_1_Z[376:0]), //o
    .io_rData_1_T (ram_io_rData_1_T[376:0]), //o
    .clk          (clk                    ), //i
    .resetn       (resetn                 )  //i
  );
  assign io_rData_0_X = _zz_io_rData_0_X;
  assign io_rData_0_Y = _zz_io_rData_0_Y;
  assign io_rData_0_Z = _zz_io_rData_0_Z;
  assign io_rData_0_T = _zz_io_rData_0_T;
  assign io_rData_1_X = _zz_io_rData_1_X;
  assign io_rData_1_Y = _zz_io_rData_1_Y;
  assign io_rData_1_Z = _zz_io_rData_1_Z;
  assign io_rData_1_T = _zz_io_rData_1_T;
  always @(posedge clk) begin
    _zz_io_rData_0_X <= (io_state_0 ? ram_io_rData_0_X : io_pInit_X);
    _zz_io_rData_0_Y <= (io_state_0 ? ram_io_rData_0_Y : io_pInit_Y);
    _zz_io_rData_0_Z <= (io_state_0 ? ram_io_rData_0_Z : io_pInit_Z);
    _zz_io_rData_0_T <= (io_state_0 ? ram_io_rData_0_T : io_pInit_T);
    _zz_io_rData_1_X <= (io_state_1 ? ram_io_rData_1_X : io_pInit_X);
    _zz_io_rData_1_Y <= (io_state_1 ? ram_io_rData_1_Y : io_pInit_Y);
    _zz_io_rData_1_Z <= (io_state_1 ? ram_io_rData_1_Z : io_pInit_Z);
    _zz_io_rData_1_T <= (io_state_1 ? ram_io_rData_1_T : io_pInit_T);
  end


endmodule

//StateRam_1 replaced by StateRam

module StateRam (
  input               io_we_0,
  input               io_we_1,
  input      [15:0]   io_address_0,
  input      [15:0]   io_address_1,
  output              io_state_0,
  output              io_state_1,
  input               io_flush,
  input      [15:0]   io_flushCnt,
  input               clk,
  input               resetn
);

  reg                 rams_0_0_io_we;
  reg        [15:0]   rams_0_0_io_wAddress;
  reg                 rams_0_0_io_wData;
  reg                 rams_0_1_io_we;
  reg        [15:0]   rams_0_1_io_wAddress;
  reg                 rams_0_1_io_wData;
  reg                 rams_1_0_io_we;
  reg        [15:0]   rams_1_0_io_wAddress;
  reg                 rams_1_0_io_wData;
  reg                 rams_1_1_io_we;
  reg        [15:0]   rams_1_1_io_wAddress;
  reg                 rams_1_1_io_wData;
  wire                rams_0_0_io_rData;
  wire                rams_0_1_io_rData;
  wire                rams_1_0_io_rData;
  wire                rams_1_1_io_rData;
  reg                 io_we_delay_1_0;
  reg                 io_we_delay_1_1;
  reg                 io_we_delay_2_0;
  reg                 io_we_delay_2_1;
  reg                 io_we_delay_3_0;
  reg                 io_we_delay_3_1;
  reg                 readArea_we_0;
  reg                 readArea_we_1;
  reg        [15:0]   io_address_regNext_0;
  reg        [15:0]   io_address_regNext_1;
  wire       [15:0]   readArea_address_0_0;
  wire       [15:0]   readArea_address_0_1;
  reg        [15:0]   readArea_address_1_0;
  reg        [15:0]   readArea_address_1_1;
  reg        [15:0]   readArea_address_2_0;
  reg        [15:0]   readArea_address_2_1;
  reg        [15:0]   readArea_address_3_0;
  reg        [15:0]   readArea_address_3_1;
  reg                 readArea_needFlip_0_0_0;
  reg                 readArea_needFlip_0_0_1;
  reg                 readArea_needFlip_0_1_0;
  reg                 readArea_needFlip_0_1_1;
  reg                 readArea_needFlip_1_0_0;
  reg                 readArea_needFlip_1_0_1;
  reg                 readArea_needFlip_1_1_0;
  reg                 readArea_needFlip_1_1_1;
  reg                 readArea_needFlip_2_0_0;
  reg                 readArea_needFlip_2_0_1;
  reg                 readArea_needFlip_2_1_0;
  reg                 readArea_needFlip_2_1_1;
  reg        [15:0]   io_address_0_regNext;
  reg        [15:0]   io_address_0_regNext_1;
  reg        [15:0]   io_address_1_regNext;
  reg        [15:0]   io_address_1_regNext_1;
  reg                 _zz_io_state_0;
  reg                 _zz_io_state_1;
  reg                 io_flush_regNext;
  reg        [15:0]   io_flushCnt_regNext;
  reg        [15:0]   io_flushCnt_regNext_1;
  reg        [15:0]   io_flushCnt_regNext_2;
  reg        [15:0]   io_flushCnt_regNext_3;

  SDPRAM_6 rams_0_0 (
    .io_we       (rams_0_0_io_we            ), //i
    .io_wAddress (rams_0_0_io_wAddress[15:0]), //i
    .io_wData    (rams_0_0_io_wData         ), //i
    .io_re       (1'b1                      ), //i
    .io_rAddress (io_address_0_regNext[15:0]), //i
    .io_rData    (rams_0_0_io_rData         ), //o
    .clk         (clk                       ), //i
    .resetn      (resetn                    )  //i
  );
  SDPRAM_6 rams_0_1 (
    .io_we       (rams_0_1_io_we            ), //i
    .io_wAddress (rams_0_1_io_wAddress[15:0]), //i
    .io_wData    (rams_0_1_io_wData         ), //i
    .io_re       (1'b1                      ), //i
    .io_rAddress (io_address_1_regNext[15:0]), //i
    .io_rData    (rams_0_1_io_rData         ), //o
    .clk         (clk                       ), //i
    .resetn      (resetn                    )  //i
  );
  SDPRAM_6 rams_1_0 (
    .io_we       (rams_1_0_io_we              ), //i
    .io_wAddress (rams_1_0_io_wAddress[15:0]  ), //i
    .io_wData    (rams_1_0_io_wData           ), //i
    .io_re       (1'b1                        ), //i
    .io_rAddress (io_address_0_regNext_1[15:0]), //i
    .io_rData    (rams_1_0_io_rData           ), //o
    .clk         (clk                         ), //i
    .resetn      (resetn                      )  //i
  );
  SDPRAM_6 rams_1_1 (
    .io_we       (rams_1_1_io_we              ), //i
    .io_wAddress (rams_1_1_io_wAddress[15:0]  ), //i
    .io_wData    (rams_1_1_io_wData           ), //i
    .io_re       (1'b1                        ), //i
    .io_rAddress (io_address_1_regNext_1[15:0]), //i
    .io_rData    (rams_1_1_io_rData           ), //o
    .clk         (clk                         ), //i
    .resetn      (resetn                      )  //i
  );
  assign readArea_address_0_0 = io_address_regNext_0;
  assign readArea_address_0_1 = io_address_regNext_1;
  assign io_state_0 = _zz_io_state_0;
  assign io_state_1 = _zz_io_state_1;
  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_0_io_wAddress = io_flushCnt_regNext;
    end else begin
      rams_0_0_io_wAddress = readArea_address_3_0;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_1_io_wAddress = io_flushCnt_regNext_1;
    end else begin
      rams_0_1_io_wAddress = readArea_address_3_0;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_0_io_wAddress = io_flushCnt_regNext_2;
    end else begin
      rams_1_0_io_wAddress = readArea_address_3_1;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_1_io_wAddress = io_flushCnt_regNext_3;
    end else begin
      rams_1_1_io_wAddress = readArea_address_3_1;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_0_io_wData = 1'b0;
    end else begin
      rams_0_0_io_wData = (! (rams_0_0_io_rData ^ readArea_needFlip_2_0_0));
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_1_io_wData = 1'b0;
    end else begin
      rams_0_1_io_wData = (! (rams_0_0_io_rData ^ readArea_needFlip_2_0_0));
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_0_io_wData = 1'b0;
    end else begin
      rams_1_0_io_wData = (! (rams_1_1_io_rData ^ readArea_needFlip_2_1_1));
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_1_io_wData = 1'b0;
    end else begin
      rams_1_1_io_wData = (! (rams_1_1_io_rData ^ readArea_needFlip_2_1_1));
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_0_io_we = 1'b1;
    end else begin
      rams_0_0_io_we = readArea_we_0;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_1_io_we = 1'b1;
    end else begin
      rams_0_1_io_we = readArea_we_0;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_0_io_we = 1'b1;
    end else begin
      rams_1_0_io_we = readArea_we_1;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_1_io_we = 1'b1;
    end else begin
      rams_1_1_io_we = readArea_we_1;
    end
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      io_we_delay_1_0 <= 1'b0;
      io_we_delay_1_1 <= 1'b0;
      io_we_delay_2_0 <= 1'b0;
      io_we_delay_2_1 <= 1'b0;
      io_we_delay_3_0 <= 1'b0;
      io_we_delay_3_1 <= 1'b0;
      readArea_we_0 <= 1'b0;
      readArea_we_1 <= 1'b0;
    end else begin
      io_we_delay_1_0 <= io_we_0;
      io_we_delay_1_1 <= io_we_1;
      io_we_delay_2_0 <= io_we_delay_1_0;
      io_we_delay_2_1 <= io_we_delay_1_1;
      io_we_delay_3_0 <= io_we_delay_2_0;
      io_we_delay_3_1 <= io_we_delay_2_1;
      readArea_we_0 <= io_we_delay_3_0;
      readArea_we_1 <= io_we_delay_3_1;
    end
  end

  always @(posedge clk) begin
    io_address_regNext_0 <= io_address_0;
    io_address_regNext_1 <= io_address_1;
    readArea_address_1_0 <= readArea_address_0_0;
    readArea_address_1_1 <= readArea_address_0_1;
    readArea_address_2_0 <= readArea_address_1_0;
    readArea_address_2_1 <= readArea_address_1_1;
    readArea_address_3_0 <= readArea_address_2_0;
    readArea_address_3_1 <= readArea_address_2_1;
    io_address_0_regNext <= io_address_0;
    io_address_0_regNext_1 <= io_address_0;
    io_address_1_regNext <= io_address_1;
    io_address_1_regNext_1 <= io_address_1;
    readArea_needFlip_0_0_0 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_0_0)) ^ 1'b0);
    readArea_needFlip_0_0_1 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_0_1)) ^ 1'b0);
    readArea_needFlip_0_1_0 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_0_0)) ^ 1'b0);
    readArea_needFlip_0_1_1 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_0_1)) ^ 1'b0);
    readArea_needFlip_1_0_0 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_1_0)) ^ readArea_needFlip_0_0_0);
    readArea_needFlip_1_0_1 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_1_1)) ^ readArea_needFlip_0_0_1);
    readArea_needFlip_1_1_0 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_1_0)) ^ readArea_needFlip_0_1_0);
    readArea_needFlip_1_1_1 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_1_1)) ^ readArea_needFlip_0_1_1);
    readArea_needFlip_2_0_0 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_2_0)) ^ readArea_needFlip_1_0_0);
    readArea_needFlip_2_0_1 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_2_1)) ^ readArea_needFlip_1_0_1);
    readArea_needFlip_2_1_0 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_2_0)) ^ readArea_needFlip_1_1_0);
    readArea_needFlip_2_1_1 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_2_1)) ^ readArea_needFlip_1_1_1);
    _zz_io_state_0 <= ((rams_0_0_io_rData ^ rams_1_0_io_rData) ^ (readArea_needFlip_2_0_0 ^ readArea_needFlip_2_1_0));
    _zz_io_state_1 <= ((rams_0_1_io_rData ^ rams_1_1_io_rData) ^ (readArea_needFlip_2_0_1 ^ readArea_needFlip_2_1_1));
    io_flush_regNext <= io_flush;
  end

  always @(posedge clk) begin
    io_flushCnt_regNext <= io_flushCnt;
    io_flushCnt_regNext_1 <= io_flushCnt;
    io_flushCnt_regNext_2 <= io_flushCnt;
    io_flushCnt_regNext_3 <= io_flushCnt;
  end


endmodule

module BADD (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  input               io_c,
  output     [377:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [56:0]   adder_adds_5_io_A_0;
  wire       [56:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [57:0]   adder_adds_5_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [63:0]   _zz_io_A_0_6;
  reg        [63:0]   _zz_io_A_0_7;
  reg        [63:0]   _zz_io_A_0_8;
  reg        [63:0]   _zz_io_A_0_9;
  reg        [56:0]   _zz_io_A_0_10;
  reg        [56:0]   _zz_io_A_0_11;
  reg        [56:0]   _zz_io_A_0_12;
  reg        [56:0]   _zz_io_A_0_13;
  reg        [56:0]   _zz_io_A_0_14;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [63:0]   _zz_io_A_1_6;
  reg        [63:0]   _zz_io_A_1_7;
  reg        [63:0]   _zz_io_A_1_8;
  reg        [63:0]   _zz_io_A_1_9;
  reg        [56:0]   _zz_io_A_1_10;
  reg        [56:0]   _zz_io_A_1_11;
  reg        [56:0]   _zz_io_A_1_12;
  reg        [56:0]   _zz_io_A_1_13;
  reg        [56:0]   _zz_io_A_1_14;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  reg        [56:0]   _zz_io_s_21;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_167 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[56:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[56:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[57:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_5_io_A_0 = _zz_io_A_0_14;
  assign adder_adds_0_io_A_1 = (~ io_b[63 : 0]);
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign adder_adds_5_io_A_1 = _zz_io_A_1_14;
  assign io_s = {_zz_io_s,{_zz_io_s_21,{_zz_io_s_20,{_zz_io_s_18,{_zz_io_s_15,{_zz_io_s_11,_zz_io_s_6}}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[319 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_0_10 <= io_a[376 : 320];
    _zz_io_A_0_11 <= _zz_io_A_0_10;
    _zz_io_A_0_12 <= _zz_io_A_0_11;
    _zz_io_A_0_13 <= _zz_io_A_0_12;
    _zz_io_A_0_14 <= _zz_io_A_0_13;
    _zz_io_A_1 <= (~ io_b[127 : 64]);
    _zz_io_A_1_1 <= (~ io_b[191 : 128]);
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= (~ io_b[255 : 192]);
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= (~ io_b[319 : 256]);
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_A_1_10 <= (~ io_b[376 : 320]);
    _zz_io_A_1_11 <= _zz_io_A_1_10;
    _zz_io_A_1_12 <= _zz_io_A_1_11;
    _zz_io_A_1_13 <= _zz_io_A_1_12;
    _zz_io_A_1_14 <= _zz_io_A_1_13;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= (! adder_adds_5_io_S[57]);
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_8 <= _zz_io_s_7;
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_21 <= adder_adds_5_io_S[56 : 0];
  end


endmodule

//FineReduction replaced by FineReduction_1

//MADD_7 replaced by MADD_12

//MADD_6 replaced by MADD_12

//MADD_5 replaced by MADD_12

//MADD_4 replaced by MADD_12

//MADD_3 replaced by MADD_8

//MADD_2 replaced by MADD_8

//MADD_1 replaced by MADD_8

//MADD replaced by MADD_8

//KaratsubaMMUL_8 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_7 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_6 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_5 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_4 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_3 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_2 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_1 replaced by KaratsubaMMUL_9

//KaratsubaMMUL replaced by KaratsubaMMUL_9

module FineReduction_1 (
  input      [377:0]  io_a,
  output     [376:0]  io_r,
  input               clk,
  input               resetn
);

  wire       [378:0]  singleAdd_add_io_s;
  wire       [376:0]  _zz__zz_io_r;
  wire       [376:0]  _zz__zz_io_r_1;
  reg        [377:0]  io_a_delay_1;
  reg        [377:0]  io_a_delay_2;
  reg        [377:0]  io_a_delay_3;
  reg        [377:0]  io_a_delay_4;
  reg        [377:0]  io_a_delay_5;
  reg        [377:0]  singleAdd_a;
  reg        [376:0]  _zz_io_r;

  assign _zz__zz_io_r = singleAdd_a[376:0];
  assign _zz__zz_io_r_1 = singleAdd_add_io_s[376:0];
  BADD_19 singleAdd_add (
    .io_a   (io_a[377:0]                                                                                         ), //i
    .io_b   (378'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001), //i
    .io_c   (1'b1                                                                                                ), //i
    .io_s   (singleAdd_add_io_s[378:0]                                                                           ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  assign io_r = _zz_io_r;
  always @(posedge clk) begin
    io_a_delay_1 <= io_a;
    io_a_delay_2 <= io_a_delay_1;
    io_a_delay_3 <= io_a_delay_2;
    io_a_delay_4 <= io_a_delay_3;
    io_a_delay_5 <= io_a_delay_4;
    singleAdd_a <= io_a_delay_5;
    _zz_io_r <= (singleAdd_add_io_s[377] ? _zz__zz_io_r : _zz__zz_io_r_1);
  end


endmodule

//MADD_15 replaced by MADD_12

//MADD_14 replaced by MADD_12

//MADD_13 replaced by MADD_12

module MADD_12 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  output     [376:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [377:0]  add_11604_io_s;
  wire       [376:0]  reduction_io_r;

  BADD_23 add_11604 (
    .io_a   (io_a[376:0]          ), //i
    .io_b   (io_b[376:0]          ), //i
    .io_c   (1'b1                 ), //i
    .io_s   (add_11604_io_s[377:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  FineReduction_53 reduction (
    .io_a   (add_11604_io_s[377:0]), //i
    .io_r   (reduction_io_r[376:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign io_s = reduction_io_r;

endmodule

//MADD_11 replaced by MADD_8

//MADD_10 replaced by MADD_8

//MADD_9 replaced by MADD_8

module MADD_8 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  output     [376:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [377:0]  add_11604_io_s;
  wire       [376:0]  reduction_io_r;

  BADD_27 add_11604 (
    .io_a   (io_a[376:0]          ), //i
    .io_b   (io_b[376:0]          ), //i
    .io_c   (1'b0                 ), //i
    .io_s   (add_11604_io_s[377:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  FineReduction_26 reduction (
    .io_a   (add_11604_io_s[377:0]), //i
    .io_r   (reduction_io_r[376:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign io_s = reduction_io_r;

endmodule

//KaratsubaMMUL_17 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_16 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_15 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_14 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_13 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_12 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_11 replaced by KaratsubaMMUL_9

//KaratsubaMMUL_10 replaced by KaratsubaMMUL_9

module KaratsubaMMUL_9 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  output     [376:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [377:0]  useBarrett_cMul1_io_a;
  wire       [377:0]  useBarrett_cMul2_io_a;
  wire       [378:0]  useBarrett_reduction_io_a;
  wire       [753:0]  useBarrett_mul_io_p;
  wire       [755:0]  useBarrett_cMul1_io_p;
  wire       [378:0]  useBarrett_cMul2_io_p;
  wire       [379:0]  useBarrett_sub_io_s;
  wire       [376:0]  useBarrett_reduction_io_r;
  reg        [378:0]  _zz_io_a;
  reg        [378:0]  _zz_io_a_1;
  reg        [378:0]  _zz_io_a_2;
  reg        [378:0]  _zz_io_a_3;
  reg        [378:0]  _zz_io_a_4;
  reg        [378:0]  _zz_io_a_5;
  reg        [378:0]  _zz_io_a_6;
  reg        [378:0]  _zz_io_a_7;
  reg        [378:0]  _zz_io_a_8;
  reg        [378:0]  _zz_io_a_9;
  reg        [378:0]  _zz_io_a_10;
  reg        [378:0]  _zz_io_a_11;
  reg        [378:0]  _zz_io_a_12;
  reg        [378:0]  _zz_io_a_13;
  reg        [378:0]  _zz_io_a_14;
  reg        [378:0]  _zz_io_a_15;
  reg        [378:0]  _zz_io_a_16;
  reg        [378:0]  _zz_io_a_17;
  reg        [378:0]  _zz_io_a_18;
  reg        [378:0]  _zz_io_a_19;
  reg        [378:0]  _zz_io_a_20;
  reg        [378:0]  _zz_io_a_21;
  reg        [378:0]  _zz_io_a_22;
  reg        [378:0]  _zz_io_a_23;
  reg        [378:0]  _zz_io_a_24;
  reg        [378:0]  _zz_io_a_25;
  reg        [378:0]  _zz_io_a_26;
  reg        [378:0]  _zz_io_a_27;
  reg        [378:0]  _zz_io_a_28;
  reg        [378:0]  _zz_io_a_29;
  reg        [378:0]  _zz_io_a_30;
  reg        [378:0]  _zz_io_a_31;
  reg        [378:0]  _zz_io_a_32;
  reg        [378:0]  _zz_io_a_33;
  reg        [378:0]  _zz_io_a_34;
  reg        [378:0]  _zz_io_a_35;
  reg        [378:0]  _zz_io_a_36;
  reg        [378:0]  _zz_io_a_37;
  reg        [378:0]  _zz_io_a_38;
  reg        [378:0]  _zz_io_a_39;
  reg        [378:0]  _zz_io_a_40;

  KaratsubaMUL_34 useBarrett_mul (
    .io_a   (io_a[376:0]               ), //i
    .io_b   (io_b[376:0]               ), //i
    .io_p   (useBarrett_mul_io_p[753:0]), //o
    .clk    (clk                       ), //i
    .resetn (resetn                    )  //i
  );
  KaratsubaMUL_35 useBarrett_cMul1 (
    .io_a   (useBarrett_cMul1_io_a[377:0]                                                                        ), //i
    .io_b   (378'h261508d0cc4060e976c3ca0582ef4f73bbad0de6776b1a06af2d488d85a6d02d0ed687789c42a591f9fd58c5e4daffc), //i
    .io_p   (useBarrett_cMul1_io_p[755:0]                                                                        ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  BCMUL_17 useBarrett_cMul2 (
    .io_a   (useBarrett_cMul2_io_a[377:0]), //i
    .io_p   (useBarrett_cMul2_io_p[378:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_36 useBarrett_sub (
    .io_a   (_zz_io_a_40[378:0]          ), //i
    .io_b   (useBarrett_cMul2_io_p[378:0]), //i
    .io_c   (1'b1                        ), //i
    .io_s   (useBarrett_sub_io_s[379:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  FineReduction_35 useBarrett_reduction (
    .io_a   (useBarrett_reduction_io_a[378:0]), //i
    .io_r   (useBarrett_reduction_io_r[376:0]), //o
    .clk    (clk                             ), //i
    .resetn (resetn                          )  //i
  );
  assign useBarrett_cMul1_io_a = useBarrett_mul_io_p[753 : 376];
  assign useBarrett_cMul2_io_a = useBarrett_cMul1_io_p[755 : 378];
  assign useBarrett_reduction_io_a = useBarrett_sub_io_s[378:0];
  assign io_p = useBarrett_reduction_io_r;
  always @(posedge clk) begin
    _zz_io_a <= useBarrett_mul_io_p[378:0];
    _zz_io_a_1 <= _zz_io_a;
    _zz_io_a_2 <= _zz_io_a_1;
    _zz_io_a_3 <= _zz_io_a_2;
    _zz_io_a_4 <= _zz_io_a_3;
    _zz_io_a_5 <= _zz_io_a_4;
    _zz_io_a_6 <= _zz_io_a_5;
    _zz_io_a_7 <= _zz_io_a_6;
    _zz_io_a_8 <= _zz_io_a_7;
    _zz_io_a_9 <= _zz_io_a_8;
    _zz_io_a_10 <= _zz_io_a_9;
    _zz_io_a_11 <= _zz_io_a_10;
    _zz_io_a_12 <= _zz_io_a_11;
    _zz_io_a_13 <= _zz_io_a_12;
    _zz_io_a_14 <= _zz_io_a_13;
    _zz_io_a_15 <= _zz_io_a_14;
    _zz_io_a_16 <= _zz_io_a_15;
    _zz_io_a_17 <= _zz_io_a_16;
    _zz_io_a_18 <= _zz_io_a_17;
    _zz_io_a_19 <= _zz_io_a_18;
    _zz_io_a_20 <= _zz_io_a_19;
    _zz_io_a_21 <= _zz_io_a_20;
    _zz_io_a_22 <= _zz_io_a_21;
    _zz_io_a_23 <= _zz_io_a_22;
    _zz_io_a_24 <= _zz_io_a_23;
    _zz_io_a_25 <= _zz_io_a_24;
    _zz_io_a_26 <= _zz_io_a_25;
    _zz_io_a_27 <= _zz_io_a_26;
    _zz_io_a_28 <= _zz_io_a_27;
    _zz_io_a_29 <= _zz_io_a_28;
    _zz_io_a_30 <= _zz_io_a_29;
    _zz_io_a_31 <= _zz_io_a_30;
    _zz_io_a_32 <= _zz_io_a_31;
    _zz_io_a_33 <= _zz_io_a_32;
    _zz_io_a_34 <= _zz_io_a_33;
    _zz_io_a_35 <= _zz_io_a_34;
    _zz_io_a_36 <= _zz_io_a_35;
    _zz_io_a_37 <= _zz_io_a_36;
    _zz_io_a_38 <= _zz_io_a_37;
    _zz_io_a_39 <= _zz_io_a_38;
    _zz_io_a_40 <= _zz_io_a_39;
  end


endmodule

//SDPRAM replaced by SDPRAM_1

module SDPRAM_1 (
  input               io_we,
  input      [7:0]    io_wAddress,
  input      [376:0]  io_wData_a_X,
  input      [376:0]  io_wData_a_Y,
  input      [376:0]  io_wData_a_Z,
  input      [376:0]  io_wData_a_T,
  input      [376:0]  io_wData_b_X,
  input      [376:0]  io_wData_b_Y,
  input      [376:0]  io_wData_b_Z,
  input      [376:0]  io_wData_b_T,
  input      [15:0]   io_wData_address,
  input               io_re,
  input      [7:0]    io_rAddress,
  output     [376:0]  io_rData_a_X,
  output     [376:0]  io_rData_a_Y,
  output     [376:0]  io_rData_a_Z,
  output     [376:0]  io_rData_a_T,
  output     [376:0]  io_rData_b_X,
  output     [376:0]  io_rData_b_Y,
  output     [376:0]  io_rData_b_Z,
  output     [376:0]  io_rData_b_T,
  output     [15:0]   io_rData_address,
  input               clk,
  input               resetn
);

  wire       [3031:0] ram_doutb;
  reg        [7:0]    io_wAddress_regNext;
  reg        [3031:0] _zz_dina;
  reg                 io_we_regNext;
  reg        [7:0]    io_rAddress_regNext;
  reg                 io_re_regNext;
  wire       [1507:0] _zz_io_rData_a_X;
  wire       [1507:0] _zz_io_rData_b_X;

  xpm_memory_sdpram #(
    .ADDR_WIDTH_A(8),
    .ADDR_WIDTH_B(8),
    .AUTO_SLEEP_TIME(0),
    .BYTE_WRITE_WIDTH_A(3032),
    .CASCADE_HEIGHT(0),
    .CLOCKING_MODE("common_clock"),
    .ECC_MODE("no_ecc"),
    .MEMORY_INIT_FILE("none"),
    .MEMORY_INIT_PARAM("0"),
    .MEMORY_OPTIMIZATION("true"),
    .MEMORY_PRIMITIVE("auto"),
    .MEMORY_SIZE(776192),
    .MESSAGE_CONTROL(0),
    .READ_DATA_WIDTH_B(3032),
    .READ_LATENCY_B(3),
    .READ_RESET_VALUE_B("0"),
    .RST_MODE_A("SYNC"),
    .RST_MODE_B("SYNC"),
    .SIM_ASSERT_CHK(0),
    .USE_EMBEDDED_CONSTRAINT(0),
    .USE_MEM_INIT(1),
    .WAKEUP_TIME("disable_sleep"),
    .WRITE_DATA_WIDTH_A(3032),
    .WRITE_MODE_B("read_first"),
    .WRITE_PROTECT(1)
  ) ram (
    .addra          (io_wAddress_regNext[7:0]), //i
    .addrb          (io_rAddress_regNext[7:0]), //i
    .dina           (_zz_dina[3031:0]        ), //i
    .doutb          (ram_doutb[3031:0]       ), //o
    .enb            (io_re_regNext           ), //i
    .wea            (io_we_regNext           ), //i
    .clka           (clk                     ), //i
    .clkb           (clk                     ), //i
    .ena            (1'b1                    ), //i
    .injectdbiterra (1'b0                    ), //i
    .injectsbiterra (1'b0                    ), //i
    .regceb         (1'b1                    ), //i
    .rstb           (1'b0                    ), //i
    .sleep          (1'b0                    )  //i
  );
  assign _zz_io_rData_a_X = ram_doutb[1507 : 0];
  assign io_rData_a_X = _zz_io_rData_a_X[376 : 0];
  assign io_rData_a_Y = _zz_io_rData_a_X[753 : 377];
  assign io_rData_a_Z = _zz_io_rData_a_X[1130 : 754];
  assign io_rData_a_T = _zz_io_rData_a_X[1507 : 1131];
  assign _zz_io_rData_b_X = ram_doutb[3015 : 1508];
  assign io_rData_b_X = _zz_io_rData_b_X[376 : 0];
  assign io_rData_b_Y = _zz_io_rData_b_X[753 : 377];
  assign io_rData_b_Z = _zz_io_rData_b_X[1130 : 754];
  assign io_rData_b_T = _zz_io_rData_b_X[1507 : 1131];
  assign io_rData_address = ram_doutb[3031 : 3016];
  always @(posedge clk) begin
    io_wAddress_regNext <= io_wAddress;
    _zz_dina <= {io_wData_address,{{io_wData_b_T,{io_wData_b_Z,{io_wData_b_Y,io_wData_b_X}}},{io_wData_a_T,{io_wData_a_Z,{io_wData_a_Y,io_wData_a_X}}}}};
    io_we_regNext <= io_we;
    io_rAddress_regNext <= io_rAddress;
    io_re_regNext <= io_re;
  end


endmodule

//TDPRAM replaced by TDPRAM_1

module TDPRAM_1 (
  input               io_we_0,
  input               io_we_1,
  input      [15:0]   io_address_0,
  input      [15:0]   io_address_1,
  input      [376:0]  io_wData_0_X,
  input      [376:0]  io_wData_0_Y,
  input      [376:0]  io_wData_0_Z,
  input      [376:0]  io_wData_0_T,
  input      [376:0]  io_wData_1_X,
  input      [376:0]  io_wData_1_Y,
  input      [376:0]  io_wData_1_Z,
  input      [376:0]  io_wData_1_T,
  input               io_ce_0,
  input               io_ce_1,
  output     [376:0]  io_rData_0_X,
  output     [376:0]  io_rData_0_Y,
  output     [376:0]  io_rData_0_Z,
  output     [376:0]  io_rData_0_T,
  output     [376:0]  io_rData_1_X,
  output     [376:0]  io_rData_1_Y,
  output     [376:0]  io_rData_1_Z,
  output     [376:0]  io_rData_1_T,
  input               clk,
  input               resetn
);

  wire       [1507:0] ram_douta;
  wire       [1507:0] ram_doutb;
  reg        [15:0]   io_address_0_regNext;
  reg        [1507:0] _zz_dina;
  reg                 io_ce_0_regNext;
  reg                 io_we_0_regNext;
  reg        [15:0]   io_address_1_regNext;
  reg        [1507:0] _zz_dinb;
  reg                 io_ce_1_regNext;
  reg                 io_we_1_regNext;

  xpm_memory_tdpram #(
    .ADDR_WIDTH_A(16),
    .ADDR_WIDTH_B(16),
    .AUTO_SLEEP_TIME(0),
    .BYTE_WRITE_WIDTH_A(1508),
    .BYTE_WRITE_WIDTH_B(1508),
    .CASCADE_HEIGHT(0),
    .CLOCKING_MODE("common_clock"),
    .ECC_MODE("no_ecc"),
    .MEMORY_INIT_FILE("none"),
    .MEMORY_INIT_PARAM("0"),
    .MEMORY_OPTIMIZATION("true"),
    .MEMORY_PRIMITIVE("ultra"),
    .MEMORY_SIZE(61767680),
    .MESSAGE_CONTROL(0),
    .READ_DATA_WIDTH_A(1508),
    .READ_DATA_WIDTH_B(1508),
    .READ_LATENCY_A(28),
    .READ_LATENCY_B(28),
    .READ_RESET_VALUE_A("0"),
    .READ_RESET_VALUE_B("0"),
    .RST_MODE_A("SYNC"),
    .RST_MODE_B("SYNC"),
    .SIM_ASSERT_CHK(0),
    .USE_EMBEDDED_CONSTRAINT(0),
    .USE_MEM_INIT(1),
    .USE_MEM_INIT_MMI(0),
    .WAKEUP_TIME("disable_sleep"),
    .WRITE_DATA_WIDTH_A(1508),
    .WRITE_DATA_WIDTH_B(1508),
    .WRITE_MODE_A("no_change"),
    .WRITE_MODE_B("no_change"),
    .WRITE_PROTECT(1)
  ) ram (
    .addra          (io_address_0_regNext[15:0]), //i
    .addrb          (io_address_1_regNext[15:0]), //i
    .dina           (_zz_dina[1507:0]          ), //i
    .dinb           (_zz_dinb[1507:0]          ), //i
    .douta          (ram_douta[1507:0]         ), //o
    .doutb          (ram_doutb[1507:0]         ), //o
    .ena            (io_ce_0_regNext           ), //i
    .enb            (io_ce_1_regNext           ), //i
    .wea            (io_we_0_regNext           ), //i
    .web            (io_we_1_regNext           ), //i
    .clka           (clk                       ), //i
    .clkb           (clk                       ), //i
    .injectdbiterra (1'b0                      ), //i
    .injectdbiterrb (1'b0                      ), //i
    .injectsbiterra (1'b0                      ), //i
    .injectsbiterrb (1'b0                      ), //i
    .regcea         (1'b1                      ), //i
    .regceb         (1'b1                      ), //i
    .rsta           (1'b0                      ), //i
    .rstb           (1'b0                      ), //i
    .sleep          (1'b0                      )  //i
  );
  assign io_rData_0_X = ram_douta[376 : 0];
  assign io_rData_0_Y = ram_douta[753 : 377];
  assign io_rData_0_Z = ram_douta[1130 : 754];
  assign io_rData_0_T = ram_douta[1507 : 1131];
  assign io_rData_1_X = ram_doutb[376 : 0];
  assign io_rData_1_Y = ram_doutb[753 : 377];
  assign io_rData_1_Z = ram_doutb[1130 : 754];
  assign io_rData_1_T = ram_doutb[1507 : 1131];
  always @(posedge clk) begin
    io_address_0_regNext <= io_address_0;
    _zz_dina <= {io_wData_0_T,{io_wData_0_Z,{io_wData_0_Y,io_wData_0_X}}};
    io_ce_0_regNext <= io_ce_0;
    io_we_0_regNext <= io_we_0;
    io_address_1_regNext <= io_address_1;
    _zz_dinb <= {io_wData_1_T,{io_wData_1_Z,{io_wData_1_Y,io_wData_1_X}}};
    io_ce_1_regNext <= io_ce_1;
    io_we_1_regNext <= io_we_1;
  end


endmodule

//SDPRAM_5 replaced by SDPRAM_6

//SDPRAM_4 replaced by SDPRAM_6

//SDPRAM_3 replaced by SDPRAM_6

//SDPRAM_2 replaced by SDPRAM_6

//SDPRAM_9 replaced by SDPRAM_6

//SDPRAM_8 replaced by SDPRAM_6

//SDPRAM_7 replaced by SDPRAM_6

module SDPRAM_6 (
  input               io_we,
  input      [15:0]   io_wAddress,
  input               io_wData,
  input               io_re,
  input      [15:0]   io_rAddress,
  output              io_rData,
  input               clk,
  input               resetn
);

  wire       [0:0]    ram_doutb;
  reg        [15:0]   io_wAddress_regNext;
  reg        [0:0]    _zz_dina;
  reg                 io_we_regNext;
  reg        [15:0]   io_rAddress_regNext;
  reg                 io_re_regNext;

  xpm_memory_sdpram #(
    .ADDR_WIDTH_A(16),
    .ADDR_WIDTH_B(16),
    .AUTO_SLEEP_TIME(0),
    .BYTE_WRITE_WIDTH_A(1),
    .CASCADE_HEIGHT(0),
    .CLOCKING_MODE("common_clock"),
    .ECC_MODE("no_ecc"),
    .MEMORY_INIT_FILE("none"),
    .MEMORY_INIT_PARAM("0"),
    .MEMORY_OPTIMIZATION("true"),
    .MEMORY_PRIMITIVE("auto"),
    .MEMORY_SIZE(40960),
    .MESSAGE_CONTROL(0),
    .READ_DATA_WIDTH_B(1),
    .READ_LATENCY_B(2),
    .READ_RESET_VALUE_B("0"),
    .RST_MODE_A("SYNC"),
    .RST_MODE_B("SYNC"),
    .SIM_ASSERT_CHK(0),
    .USE_EMBEDDED_CONSTRAINT(0),
    .USE_MEM_INIT(1),
    .WAKEUP_TIME("disable_sleep"),
    .WRITE_DATA_WIDTH_A(1),
    .WRITE_MODE_B("read_first"),
    .WRITE_PROTECT(1)
  ) ram (
    .addra          (io_wAddress_regNext[15:0]), //i
    .addrb          (io_rAddress_regNext[15:0]), //i
    .dina           (_zz_dina                 ), //i
    .doutb          (ram_doutb                ), //o
    .enb            (io_re_regNext            ), //i
    .wea            (io_we_regNext            ), //i
    .clka           (clk                      ), //i
    .clkb           (clk                      ), //i
    .ena            (1'b1                     ), //i
    .injectdbiterra (1'b0                     ), //i
    .injectsbiterra (1'b0                     ), //i
    .regceb         (1'b1                     ), //i
    .rstb           (1'b0                     ), //i
    .sleep          (1'b0                     )  //i
  );
  assign io_rData = ram_doutb[0];
  always @(posedge clk) begin
    io_wAddress_regNext <= io_wAddress;
    _zz_dina <= io_wData;
    io_we_regNext <= io_we;
    io_rAddress_regNext <= io_rAddress;
    io_re_regNext <= io_re;
  end


endmodule

//ADD_5 replaced by ADD_167

//ADD_4 replaced by ADD_5756

//ADD_3 replaced by ADD_5756

//ADD_2 replaced by ADD_5756

//ADD_1 replaced by ADD_5756

//ADD replaced by ADD_5756

//BADD_1 replaced by BADD_19

//FineReduction_2 replaced by FineReduction_53

//BADD_2 replaced by BADD_23

//FineReduction_3 replaced by FineReduction_53

//BADD_3 replaced by BADD_23

//FineReduction_4 replaced by FineReduction_53

//BADD_4 replaced by BADD_23

//FineReduction_5 replaced by FineReduction_53

//BADD_5 replaced by BADD_23

//FineReduction_6 replaced by FineReduction_26

//BADD_6 replaced by BADD_27

//FineReduction_7 replaced by FineReduction_26

//BADD_7 replaced by BADD_27

//FineReduction_8 replaced by FineReduction_26

//BADD_8 replaced by BADD_27

//FineReduction_9 replaced by FineReduction_26

//BADD_9 replaced by BADD_27

//FineReduction_10 replaced by FineReduction_35

//BADD_10 replaced by BADD_36

//BCMUL replaced by BCMUL_17

//KaratsubaMUL_1 replaced by KaratsubaMUL_35

//KaratsubaMUL replaced by KaratsubaMUL_34

//FineReduction_11 replaced by FineReduction_35

//BADD_11 replaced by BADD_36

//BCMUL_1 replaced by BCMUL_17

//KaratsubaMUL_3 replaced by KaratsubaMUL_35

//KaratsubaMUL_2 replaced by KaratsubaMUL_34

//FineReduction_12 replaced by FineReduction_35

//BADD_12 replaced by BADD_36

//BCMUL_2 replaced by BCMUL_17

//KaratsubaMUL_5 replaced by KaratsubaMUL_35

//KaratsubaMUL_4 replaced by KaratsubaMUL_34

//FineReduction_13 replaced by FineReduction_35

//BADD_13 replaced by BADD_36

//BCMUL_3 replaced by BCMUL_17

//KaratsubaMUL_7 replaced by KaratsubaMUL_35

//KaratsubaMUL_6 replaced by KaratsubaMUL_34

//FineReduction_14 replaced by FineReduction_35

//BADD_14 replaced by BADD_36

//BCMUL_4 replaced by BCMUL_17

//KaratsubaMUL_9 replaced by KaratsubaMUL_35

//KaratsubaMUL_8 replaced by KaratsubaMUL_34

//FineReduction_15 replaced by FineReduction_35

//BADD_15 replaced by BADD_36

//BCMUL_5 replaced by BCMUL_17

//KaratsubaMUL_11 replaced by KaratsubaMUL_35

//KaratsubaMUL_10 replaced by KaratsubaMUL_34

//FineReduction_16 replaced by FineReduction_35

//BADD_16 replaced by BADD_36

//BCMUL_6 replaced by BCMUL_17

//KaratsubaMUL_13 replaced by KaratsubaMUL_35

//KaratsubaMUL_12 replaced by KaratsubaMUL_34

//FineReduction_17 replaced by FineReduction_35

//BADD_17 replaced by BADD_36

//BCMUL_7 replaced by BCMUL_17

//KaratsubaMUL_15 replaced by KaratsubaMUL_35

//KaratsubaMUL_14 replaced by KaratsubaMUL_34

//FineReduction_18 replaced by FineReduction_35

//BADD_18 replaced by BADD_36

//BCMUL_8 replaced by BCMUL_17

//KaratsubaMUL_17 replaced by KaratsubaMUL_35

//KaratsubaMUL_16 replaced by KaratsubaMUL_34

module BADD_19 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  input               io_c,
  output     [378:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [57:0]   adder_adds_5_io_A_0;
  wire       [57:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [58:0]   adder_adds_5_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [63:0]   _zz_io_A_0_6;
  reg        [63:0]   _zz_io_A_0_7;
  reg        [63:0]   _zz_io_A_0_8;
  reg        [63:0]   _zz_io_A_0_9;
  reg        [57:0]   _zz_io_A_0_10;
  reg        [57:0]   _zz_io_A_0_11;
  reg        [57:0]   _zz_io_A_0_12;
  reg        [57:0]   _zz_io_A_0_13;
  reg        [57:0]   _zz_io_A_0_14;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [63:0]   _zz_io_A_1_6;
  reg        [63:0]   _zz_io_A_1_7;
  reg        [63:0]   _zz_io_A_1_8;
  reg        [63:0]   _zz_io_A_1_9;
  reg        [57:0]   _zz_io_A_1_10;
  reg        [57:0]   _zz_io_A_1_11;
  reg        [57:0]   _zz_io_A_1_12;
  reg        [57:0]   _zz_io_A_1_13;
  reg        [57:0]   _zz_io_A_1_14;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  reg        [57:0]   _zz_io_s_21;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_5761 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[57:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[57:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[58:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_5_io_A_0 = _zz_io_A_0_14;
  assign adder_adds_0_io_A_1 = (~ io_b[63 : 0]);
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign adder_adds_5_io_A_1 = _zz_io_A_1_14;
  assign io_s = {_zz_io_s,{_zz_io_s_21,{_zz_io_s_20,{_zz_io_s_18,{_zz_io_s_15,{_zz_io_s_11,_zz_io_s_6}}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[319 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_0_10 <= io_a[377 : 320];
    _zz_io_A_0_11 <= _zz_io_A_0_10;
    _zz_io_A_0_12 <= _zz_io_A_0_11;
    _zz_io_A_0_13 <= _zz_io_A_0_12;
    _zz_io_A_0_14 <= _zz_io_A_0_13;
    _zz_io_A_1 <= (~ io_b[127 : 64]);
    _zz_io_A_1_1 <= (~ io_b[191 : 128]);
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= (~ io_b[255 : 192]);
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= (~ io_b[319 : 256]);
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_A_1_10 <= (~ io_b[377 : 320]);
    _zz_io_A_1_11 <= _zz_io_A_1_10;
    _zz_io_A_1_12 <= _zz_io_A_1_11;
    _zz_io_A_1_13 <= _zz_io_A_1_12;
    _zz_io_A_1_14 <= _zz_io_A_1_13;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= (! adder_adds_5_io_S[58]);
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_8 <= _zz_io_s_7;
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_21 <= adder_adds_5_io_S[57 : 0];
  end


endmodule

//FineReduction_19 replaced by FineReduction_53

//BADD_20 replaced by BADD_23

//FineReduction_20 replaced by FineReduction_53

//BADD_21 replaced by BADD_23

//FineReduction_21 replaced by FineReduction_53

//BADD_22 replaced by BADD_23

//FineReduction_22 replaced by FineReduction_53

module BADD_23 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  input               io_c,
  output     [377:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [56:0]   adder_adds_5_io_A_0;
  wire       [56:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [57:0]   adder_adds_5_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [63:0]   _zz_io_A_0_6;
  reg        [63:0]   _zz_io_A_0_7;
  reg        [63:0]   _zz_io_A_0_8;
  reg        [63:0]   _zz_io_A_0_9;
  reg        [56:0]   _zz_io_A_0_10;
  reg        [56:0]   _zz_io_A_0_11;
  reg        [56:0]   _zz_io_A_0_12;
  reg        [56:0]   _zz_io_A_0_13;
  reg        [56:0]   _zz_io_A_0_14;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [63:0]   _zz_io_A_1_6;
  reg        [63:0]   _zz_io_A_1_7;
  reg        [63:0]   _zz_io_A_1_8;
  reg        [63:0]   _zz_io_A_1_9;
  reg        [56:0]   _zz_io_A_1_10;
  reg        [56:0]   _zz_io_A_1_11;
  reg        [56:0]   _zz_io_A_1_12;
  reg        [56:0]   _zz_io_A_1_13;
  reg        [56:0]   _zz_io_A_1_14;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [56:0]   _zz_io_s_6;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_167 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[56:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[56:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[57:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_5_io_A_0 = _zz_io_A_0_14;
  assign adder_adds_0_io_A_1 = (~ io_b[63 : 0]);
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign adder_adds_5_io_A_1 = _zz_io_A_1_14;
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[319 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_0_10 <= io_a[376 : 320];
    _zz_io_A_0_11 <= _zz_io_A_0_10;
    _zz_io_A_0_12 <= _zz_io_A_0_11;
    _zz_io_A_0_13 <= _zz_io_A_0_12;
    _zz_io_A_0_14 <= _zz_io_A_0_13;
    _zz_io_A_1 <= (~ io_b[127 : 64]);
    _zz_io_A_1_1 <= (~ io_b[191 : 128]);
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= (~ io_b[255 : 192]);
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= (~ io_b[319 : 256]);
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_A_1_10 <= (~ io_b[376 : 320]);
    _zz_io_A_1_11 <= _zz_io_A_1_10;
    _zz_io_A_1_12 <= _zz_io_A_1_11;
    _zz_io_A_1_13 <= _zz_io_A_1_12;
    _zz_io_A_1_14 <= _zz_io_A_1_13;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= (! adder_adds_5_io_S[57]);
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[56 : 0];
  end


endmodule

//FineReduction_23 replaced by FineReduction_26

//BADD_24 replaced by BADD_27

//FineReduction_24 replaced by FineReduction_26

//BADD_25 replaced by BADD_27

//FineReduction_25 replaced by FineReduction_26

//BADD_26 replaced by BADD_27

module FineReduction_26 (
  input      [377:0]  io_a,
  output     [376:0]  io_r,
  input               clk,
  input               resetn
);

  wire       [378:0]  singleAdd_add_io_s;
  wire       [376:0]  _zz__zz_io_r;
  wire       [376:0]  _zz__zz_io_r_1;
  reg        [63:0]   _zz_singleAdd_a;
  reg        [63:0]   _zz_singleAdd_a_1;
  reg        [63:0]   _zz_singleAdd_a_2;
  reg        [63:0]   _zz_singleAdd_a_3;
  reg        [63:0]   _zz_singleAdd_a_4;
  reg        [63:0]   _zz_singleAdd_a_5;
  reg        [63:0]   _zz_singleAdd_a_6;
  reg        [63:0]   _zz_singleAdd_a_7;
  reg        [63:0]   _zz_singleAdd_a_8;
  reg        [63:0]   _zz_singleAdd_a_9;
  reg        [63:0]   _zz_singleAdd_a_10;
  reg        [63:0]   _zz_singleAdd_a_11;
  reg        [63:0]   _zz_singleAdd_a_12;
  reg        [63:0]   _zz_singleAdd_a_13;
  reg        [63:0]   _zz_singleAdd_a_14;
  reg        [63:0]   _zz_singleAdd_a_15;
  reg        [63:0]   _zz_singleAdd_a_16;
  reg        [63:0]   _zz_singleAdd_a_17;
  reg        [63:0]   _zz_singleAdd_a_18;
  reg        [63:0]   _zz_singleAdd_a_19;
  reg        [57:0]   _zz_singleAdd_a_20;
  wire       [377:0]  singleAdd_a;
  reg        [376:0]  _zz_io_r;

  assign _zz__zz_io_r = singleAdd_a[376:0];
  assign _zz__zz_io_r_1 = singleAdd_add_io_s[376:0];
  BADD_619 singleAdd_add (
    .io_a   (io_a[377:0]                                                                                         ), //i
    .io_b   (378'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001), //i
    .io_c   (1'b1                                                                                                ), //i
    .io_s   (singleAdd_add_io_s[378:0]                                                                           ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  assign singleAdd_a = {_zz_singleAdd_a_20,{_zz_singleAdd_a_19,{_zz_singleAdd_a_17,{_zz_singleAdd_a_14,{_zz_singleAdd_a_10,_zz_singleAdd_a_5}}}}};
  assign io_r = _zz_io_r;
  always @(posedge clk) begin
    _zz_singleAdd_a <= io_a[63 : 0];
    _zz_singleAdd_a_1 <= _zz_singleAdd_a;
    _zz_singleAdd_a_2 <= _zz_singleAdd_a_1;
    _zz_singleAdd_a_3 <= _zz_singleAdd_a_2;
    _zz_singleAdd_a_4 <= _zz_singleAdd_a_3;
    _zz_singleAdd_a_5 <= _zz_singleAdd_a_4;
    _zz_singleAdd_a_6 <= io_a[127 : 64];
    _zz_singleAdd_a_7 <= _zz_singleAdd_a_6;
    _zz_singleAdd_a_8 <= _zz_singleAdd_a_7;
    _zz_singleAdd_a_9 <= _zz_singleAdd_a_8;
    _zz_singleAdd_a_10 <= _zz_singleAdd_a_9;
    _zz_singleAdd_a_11 <= io_a[191 : 128];
    _zz_singleAdd_a_12 <= _zz_singleAdd_a_11;
    _zz_singleAdd_a_13 <= _zz_singleAdd_a_12;
    _zz_singleAdd_a_14 <= _zz_singleAdd_a_13;
    _zz_singleAdd_a_15 <= io_a[255 : 192];
    _zz_singleAdd_a_16 <= _zz_singleAdd_a_15;
    _zz_singleAdd_a_17 <= _zz_singleAdd_a_16;
    _zz_singleAdd_a_18 <= io_a[319 : 256];
    _zz_singleAdd_a_19 <= _zz_singleAdd_a_18;
    _zz_singleAdd_a_20 <= io_a[377 : 320];
    _zz_io_r <= (singleAdd_add_io_s[377] ? _zz__zz_io_r : _zz__zz_io_r_1);
  end


endmodule

module BADD_27 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  input               io_c,
  output     [377:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [56:0]   adder_adds_5_io_A_0;
  wire       [56:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [57:0]   adder_adds_5_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [63:0]   _zz_io_A_0_6;
  reg        [63:0]   _zz_io_A_0_7;
  reg        [63:0]   _zz_io_A_0_8;
  reg        [63:0]   _zz_io_A_0_9;
  reg        [56:0]   _zz_io_A_0_10;
  reg        [56:0]   _zz_io_A_0_11;
  reg        [56:0]   _zz_io_A_0_12;
  reg        [56:0]   _zz_io_A_0_13;
  reg        [56:0]   _zz_io_A_0_14;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [63:0]   _zz_io_A_1_6;
  reg        [63:0]   _zz_io_A_1_7;
  reg        [63:0]   _zz_io_A_1_8;
  reg        [63:0]   _zz_io_A_1_9;
  reg        [56:0]   _zz_io_A_1_10;
  reg        [56:0]   _zz_io_A_1_11;
  reg        [56:0]   _zz_io_A_1_12;
  reg        [56:0]   _zz_io_A_1_13;
  reg        [56:0]   _zz_io_A_1_14;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [56:0]   _zz_io_s_6;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_167 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[56:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[56:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[57:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_5_io_A_0 = _zz_io_A_0_14;
  assign adder_adds_0_io_A_1 = io_b[63 : 0];
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign adder_adds_5_io_A_1 = _zz_io_A_1_14;
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[319 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_0_10 <= io_a[376 : 320];
    _zz_io_A_0_11 <= _zz_io_A_0_10;
    _zz_io_A_0_12 <= _zz_io_A_0_11;
    _zz_io_A_0_13 <= _zz_io_A_0_12;
    _zz_io_A_0_14 <= _zz_io_A_0_13;
    _zz_io_A_1 <= io_b[127 : 64];
    _zz_io_A_1_1 <= io_b[191 : 128];
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= io_b[255 : 192];
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= io_b[319 : 256];
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_A_1_10 <= io_b[376 : 320];
    _zz_io_A_1_11 <= _zz_io_A_1_10;
    _zz_io_A_1_12 <= _zz_io_A_1_11;
    _zz_io_A_1_13 <= _zz_io_A_1_12;
    _zz_io_A_1_14 <= _zz_io_A_1_13;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= adder_adds_5_io_S[57];
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[56 : 0];
  end


endmodule

//FineReduction_27 replaced by FineReduction_35

//BADD_28 replaced by BADD_36

//BCMUL_9 replaced by BCMUL_17

//KaratsubaMUL_19 replaced by KaratsubaMUL_35

//KaratsubaMUL_18 replaced by KaratsubaMUL_34

//FineReduction_28 replaced by FineReduction_35

//BADD_29 replaced by BADD_36

//BCMUL_10 replaced by BCMUL_17

//KaratsubaMUL_21 replaced by KaratsubaMUL_35

//KaratsubaMUL_20 replaced by KaratsubaMUL_34

//FineReduction_29 replaced by FineReduction_35

//BADD_30 replaced by BADD_36

//BCMUL_11 replaced by BCMUL_17

//KaratsubaMUL_23 replaced by KaratsubaMUL_35

//KaratsubaMUL_22 replaced by KaratsubaMUL_34

//FineReduction_30 replaced by FineReduction_35

//BADD_31 replaced by BADD_36

//BCMUL_12 replaced by BCMUL_17

//KaratsubaMUL_25 replaced by KaratsubaMUL_35

//KaratsubaMUL_24 replaced by KaratsubaMUL_34

//FineReduction_31 replaced by FineReduction_35

//BADD_32 replaced by BADD_36

//BCMUL_13 replaced by BCMUL_17

//KaratsubaMUL_27 replaced by KaratsubaMUL_35

//KaratsubaMUL_26 replaced by KaratsubaMUL_34

//FineReduction_32 replaced by FineReduction_35

//BADD_33 replaced by BADD_36

//BCMUL_14 replaced by BCMUL_17

//KaratsubaMUL_29 replaced by KaratsubaMUL_35

//KaratsubaMUL_28 replaced by KaratsubaMUL_34

//FineReduction_33 replaced by FineReduction_35

//BADD_34 replaced by BADD_36

//BCMUL_15 replaced by BCMUL_17

//KaratsubaMUL_31 replaced by KaratsubaMUL_35

//KaratsubaMUL_30 replaced by KaratsubaMUL_34

//FineReduction_34 replaced by FineReduction_35

//BADD_35 replaced by BADD_36

//BCMUL_16 replaced by BCMUL_17

//KaratsubaMUL_33 replaced by KaratsubaMUL_35

//KaratsubaMUL_32 replaced by KaratsubaMUL_34

module FineReduction_35 (
  input      [378:0]  io_a,
  output     [376:0]  io_r,
  input               clk,
  input               resetn
);

  wire       [377:0]  doubleAdd_reduction_io_a;
  wire       [378:0]  doubleAdd_add_io_s;
  wire       [376:0]  doubleAdd_reduction_io_r;
  wire       [376:0]  _zz_doubleAdd_subRom_1;
  wire       [376:0]  _zz_doubleAdd_subRom_2;
  wire       [377:0]  _zz_doubleAdd_subRom_3;
  wire       [377:0]  _zz_doubleAdd_subRom_4;
  wire       [376:0]  _zz_doubleAdd_subRom_5;
  reg        [377:0]  _zz__zz_io_b;
  wire       [2:0]    _zz__zz_io_b_1;
  wire       [377:0]  doubleAdd_subRom_0;
  wire       [377:0]  doubleAdd_subRom_1;
  wire       [377:0]  doubleAdd_subRom_2;
  wire       [377:0]  doubleAdd_subRom_3;
  wire       [377:0]  doubleAdd_subRom_4;
  wire       [377:0]  doubleAdd_subRom_5;
  wire       [377:0]  doubleAdd_subRom_6;
  wire       [377:0]  doubleAdd_subRom_7;
  reg        [377:0]  _zz_io_a;
  reg        [377:0]  _zz_io_b;

  assign _zz_doubleAdd_subRom_1 = 377'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001;
  assign _zz_doubleAdd_subRom_2 = 377'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001;
  assign _zz_doubleAdd_subRom_3 = 378'h35c748c2f8a21d58c760b80d94292763445b3e601ea271e3de6c45f741290002e16ba88600000010a11800000000002;
  assign _zz_doubleAdd_subRom_4 = 378'h35c748c2f8a21d58c760b80d94292763445b3e601ea271e3de6c45f741290002e16ba88600000010a11800000000002;
  assign _zz_doubleAdd_subRom_5 = 377'h10aaed2474f32c052b1114145e3dbb14e688dd902df3aad5cda268f2e1bd800452217cc900000018f1a400000000003;
  assign _zz__zz_io_b_1 = io_a[378 : 376];
  BADD_1124 doubleAdd_add (
    .io_a   (_zz_io_a[377:0]          ), //i
    .io_b   (_zz_io_b[377:0]          ), //i
    .io_c   (1'b1                     ), //i
    .io_s   (doubleAdd_add_io_s[378:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  FineReduction_53 doubleAdd_reduction (
    .io_a   (doubleAdd_reduction_io_a[377:0]), //i
    .io_r   (doubleAdd_reduction_io_r[376:0]), //o
    .clk    (clk                            ), //i
    .resetn (resetn                         )  //i
  );
  always @(*) begin
    case(_zz__zz_io_b_1)
      3'b000 : _zz__zz_io_b = doubleAdd_subRom_0;
      3'b001 : _zz__zz_io_b = doubleAdd_subRom_1;
      3'b010 : _zz__zz_io_b = doubleAdd_subRom_2;
      3'b011 : _zz__zz_io_b = doubleAdd_subRom_3;
      3'b100 : _zz__zz_io_b = doubleAdd_subRom_4;
      3'b101 : _zz__zz_io_b = doubleAdd_subRom_5;
      3'b110 : _zz__zz_io_b = doubleAdd_subRom_6;
      default : _zz__zz_io_b = doubleAdd_subRom_7;
    endcase
  end

  assign doubleAdd_subRom_0 = 378'h0;
  assign doubleAdd_subRom_1 = {1'd0, _zz_doubleAdd_subRom_1};
  assign doubleAdd_subRom_2 = {1'd0, _zz_doubleAdd_subRom_2};
  assign doubleAdd_subRom_3 = _zz_doubleAdd_subRom_3;
  assign doubleAdd_subRom_4 = _zz_doubleAdd_subRom_4;
  assign doubleAdd_subRom_5 = {1'd0, _zz_doubleAdd_subRom_5};
  assign doubleAdd_subRom_6 = 378'h0;
  assign doubleAdd_subRom_7 = 378'h0;
  assign doubleAdd_reduction_io_a = doubleAdd_add_io_s[377:0];
  assign io_r = doubleAdd_reduction_io_r;
  always @(posedge clk) begin
    _zz_io_a <= io_a[377:0];
    _zz_io_b <= _zz__zz_io_b;
  end


endmodule

module BADD_36 (
  input      [378:0]  io_a,
  input      [378:0]  io_b,
  input               io_c,
  output     [379:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [58:0]   adder_adds_5_io_A_0;
  wire       [58:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [59:0]   adder_adds_5_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [63:0]   _zz_io_A_0_6;
  reg        [63:0]   _zz_io_A_0_7;
  reg        [63:0]   _zz_io_A_0_8;
  reg        [63:0]   _zz_io_A_0_9;
  reg        [58:0]   _zz_io_A_0_10;
  reg        [58:0]   _zz_io_A_0_11;
  reg        [58:0]   _zz_io_A_0_12;
  reg        [58:0]   _zz_io_A_0_13;
  reg        [58:0]   _zz_io_A_0_14;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [63:0]   _zz_io_A_1_6;
  reg        [63:0]   _zz_io_A_1_7;
  reg        [63:0]   _zz_io_A_1_8;
  reg        [63:0]   _zz_io_A_1_9;
  reg        [58:0]   _zz_io_A_1_10;
  reg        [58:0]   _zz_io_A_1_11;
  reg        [58:0]   _zz_io_A_1_12;
  reg        [58:0]   _zz_io_A_1_13;
  reg        [58:0]   _zz_io_A_1_14;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  reg        [58:0]   _zz_io_s_21;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_5_io_A_0 = _zz_io_A_0_14;
  assign adder_adds_0_io_A_1 = (~ io_b[63 : 0]);
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign adder_adds_5_io_A_1 = _zz_io_A_1_14;
  assign io_s = {_zz_io_s,{_zz_io_s_21,{_zz_io_s_20,{_zz_io_s_18,{_zz_io_s_15,{_zz_io_s_11,_zz_io_s_6}}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[319 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_0_10 <= io_a[378 : 320];
    _zz_io_A_0_11 <= _zz_io_A_0_10;
    _zz_io_A_0_12 <= _zz_io_A_0_11;
    _zz_io_A_0_13 <= _zz_io_A_0_12;
    _zz_io_A_0_14 <= _zz_io_A_0_13;
    _zz_io_A_1 <= (~ io_b[127 : 64]);
    _zz_io_A_1_1 <= (~ io_b[191 : 128]);
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= (~ io_b[255 : 192]);
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= (~ io_b[319 : 256]);
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_A_1_10 <= (~ io_b[378 : 320]);
    _zz_io_A_1_11 <= _zz_io_A_1_10;
    _zz_io_A_1_12 <= _zz_io_A_1_11;
    _zz_io_A_1_13 <= _zz_io_A_1_12;
    _zz_io_A_1_14 <= _zz_io_A_1_13;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= (! adder_adds_5_io_S[59]);
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_8 <= _zz_io_s_7;
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_21 <= adder_adds_5_io_S[58 : 0];
  end


endmodule

module BCMUL_17 (
  input      [377:0]  io_a,
  output     [378:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [322:0]  NAFElements_adds_0_io_a;
  wire       [322:0]  NAFElements_adds_0_io_b;
  wire       [332:0]  NAFElements_adds_1_io_a;
  wire       [332:0]  NAFElements_adds_1_io_b;
  wire       [272:0]  NAFElements_adds_2_io_a;
  wire       [272:0]  NAFElements_adds_2_io_b;
  wire       [189:0]  NAFElements_adds_3_io_a;
  wire       [189:0]  NAFElements_adds_3_io_b;
  wire       [327:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [280:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [315:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [253:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [234:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [209:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [170:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [176:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [214:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [116:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [136:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [106:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [91:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [101:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [111:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [50:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [25:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [15:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [20:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [31:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [4:0]    adder_posMUL_multiElements_add_add_io_a;
  wire       [267:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [225:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [258:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [194:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [200:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [220:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [182:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [150:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [166:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [141:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [125:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [129:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [145:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [74:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [84:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [63:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [54:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [58:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [68:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [120:0]  adder_negMUL_multiElements_add_add_io_a;
  wire       [378:0]  adder_add_io_b;
  wire       [323:0]  NAFElements_adds_0_io_s;
  wire       [333:0]  NAFElements_adds_1_io_s;
  wire       [273:0]  NAFElements_adds_2_io_s;
  wire       [190:0]  NAFElements_adds_3_io_s;
  wire       [333:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [323:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [328:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [287:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [277:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [281:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [316:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [254:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [235:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [240:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [210:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [171:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [177:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [215:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [263:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [155:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [117:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [137:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [107:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [92:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [102:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [112:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [51:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [43:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [47:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [26:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [16:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [21:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [32:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [80:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [163:0]  adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [5:0]    adder_posMUL_multiElements_add_add_io_s;
  wire       [268:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [226:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [259:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [206:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [195:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [201:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [221:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [183:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [151:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [167:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [142:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [126:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [130:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [146:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [190:0]  adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [97:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [75:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [85:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [64:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [55:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [59:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [69:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [10:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [37:0]   adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [121:0]  adder_negMUL_multiElements_add_add_io_s;
  wire       [379:0]  adder_add_io_s;
  wire       [379:0]  _zz_io_a_11;
  wire       [378:0]  _zz_io_a_12;
  wire       [380:0]  _zz_io_a_13;
  wire       [380:0]  _zz_io_a_14;
  wire       [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  wire       [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  wire       [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  wire       [12:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  wire       [12:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  wire       [12:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  wire       [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  wire       [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  wire       [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  wire       [0:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  wire       [0:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  wire       [0:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  wire       [50:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [46:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [42:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [31:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [25:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [20:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [15:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [4:0]    _zz__zz_adder_posMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [58:0]   _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [54:0]   _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [36:0]   _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [9:0]    _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [378:0]  _zz_io_p;
  wire       [379:0]  _zz_io_p_1;
  wire       [378:0]  _zz_NAFElements_sums_0;
  reg        [63:0]   _zz_NAFElements_sums_0_1;
  reg        [63:0]   _zz_NAFElements_sums_0_2;
  reg        [63:0]   _zz_NAFElements_sums_0_3;
  reg        [63:0]   _zz_NAFElements_sums_0_4;
  reg        [63:0]   _zz_NAFElements_sums_0_5;
  reg        [63:0]   _zz_NAFElements_sums_0_6;
  reg        [63:0]   _zz_NAFElements_sums_0_7;
  reg        [63:0]   _zz_NAFElements_sums_0_8;
  reg        [63:0]   _zz_NAFElements_sums_0_9;
  reg        [63:0]   _zz_NAFElements_sums_0_10;
  reg        [58:0]   _zz_NAFElements_sums_0_11;
  reg        [58:0]   _zz_NAFElements_sums_0_12;
  reg        [58:0]   _zz_NAFElements_sums_0_13;
  reg        [58:0]   _zz_NAFElements_sums_0_14;
  reg        [58:0]   _zz_NAFElements_sums_0_15;
  wire       [378:0]  NAFElements_sums_0;
  wire       [322:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [332:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [272:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [189:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [378:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [332:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [332:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [332:0]  _zz_io_a;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [327:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [327:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [327:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  wire       [322:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [322:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [322:0]  _zz_io_a_1;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [315:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [315:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [315:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [315:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  wire       [59:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [58:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  wire       [286:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [286:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [286:0]  _zz_io_a_2;
  reg        [28:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [28:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [280:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [280:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [280:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [29:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [29:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [29:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [29:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [24:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  wire       [276:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [276:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [276:0]  _zz_io_a_3;
  reg        [3:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [3:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [34:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [262:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [11:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [11:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [11:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [11:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [6:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  wire       [253:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [253:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  wire       [61:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [2:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [2:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [2:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [58:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [58:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [2:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [8:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [239:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [239:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [239:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20;
  wire       [234:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [234:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [239:0]  _zz_io_a_4;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [214:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [214:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [214:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [214:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20;
  wire       [209:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [209:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20;
  reg        [209:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [176:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [176:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [176:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [48:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [48:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [48:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  wire       [170:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [170:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [115:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [162:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [34:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [34:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [34:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  wire       [154:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [154:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [26:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [26:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [26:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [154:0]  _zz_io_a_5;
  reg        [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [136:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [136:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [136:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [8:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [8:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [8:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  wire       [116:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [116:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [57:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [57:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [57:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [57:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [19:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [111:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [111:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [111:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [111:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  wire       [106:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [106:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [106:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [101:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [101:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [101:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  wire       [91:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [91:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [91:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [79:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  wire       [50:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [28:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [46:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [46:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [42:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [42:0]   _zz_io_a_6;
  reg        [3:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [3:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [46:0]   _zz_io_a_7;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [31:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [31:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [31:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  wire       [25:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [20:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [20:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [15:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [82:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [215:0]  _zz_adder_posMUL_multiElements_lsbMUL_p;
  wire       [4:0]    adder_posMUL_multiElements_msbMUL_p;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p_1;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p_2;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p_3;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p_4;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_1;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_2;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_3;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_4;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_5;
  reg        [373:0]  _zz_adder_posMUL_p;
  reg        [272:0]  adder_negMUL_p;
  reg        [272:0]  adder_negMUL_multiElements_lsbMUL_p;
  reg        [272:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [272:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [272:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [272:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [272:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [21:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [21:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [21:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [21:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  wire       [267:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [267:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [11:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [4:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [258:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [258:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [258:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  wire       [225:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [225:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20;
  reg        [32:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [220:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [220:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [220:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [220:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [28:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  reg        [28:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20;
  wire       [205:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [205:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20;
  reg        [205:0]  _zz_io_a_8;
  reg        [14:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [14:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [200:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [200:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [200:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [8:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  reg        [8:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20;
  wire       [194:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [194:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20;
  reg        [194:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
  reg        [5:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [51:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [189:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  wire       [61:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  wire       [182:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [182:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [54:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [54:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [54:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [166:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [166:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [166:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  wire       [150:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [150:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [15:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [166:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [145:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [145:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [145:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [145:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [17:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [17:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [17:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  wire       [141:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [141:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [129:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [129:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [129:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [1:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [1:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [1:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  wire       [125:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [125:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [61:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [15:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [82:0]   _zz_adder_negMUL_multiElements_lsbMUL_p;
  reg        [120:0]  adder_negMUL_multiElements_msbMUL_p;
  reg        [120:0]  adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [120:0]  adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [120:0]  adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [120:0]  adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [120:0]  _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [61:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [61:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [61:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [61:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [56:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [56:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [56:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [56:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  wire       [96:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [96:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [32:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [32:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [32:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [32:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [96:0]   _zz_io_a_9;
  reg        [23:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [23:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [84:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [84:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [84:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [20:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [20:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [20:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [20:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  wire       [74:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [74:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [15:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [15:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [15:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [15:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [10:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [10:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [10:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [10:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [35:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [68:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [68:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [68:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [68:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  wire       [63:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [58:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [58:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [54:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [54:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
  reg        [3:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [51:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [9:0]    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [9:0]    _zz_io_a_10;
  reg        [26:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [26:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
  reg        [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_2;
  reg        [83:0]   _zz_adder_negMUL_multiElements_msbMUL_p;
  reg        [151:0]  _zz_adder_negMUL_p;
  reg        [272:0]  adder_negMUL_p_delay_1;

  assign _zz_io_a_11 = ({2'd0,io_a} <<< 2);
  assign _zz_io_a_12 = ({1'd0,io_a} <<< 1);
  assign _zz_io_a_13 = ({3'd0,io_a} <<< 3);
  assign _zz_io_a_14 = ({3'd0,io_a} <<< 3);
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_sums_0[50:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[46:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[42:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[31:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[25:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[20:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[15:0];
  assign _zz__zz_adder_posMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[58:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_sums_0[54:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[36:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[9:0];
  assign _zz_io_p_1 = adder_add_io_s;
  assign _zz_io_p = _zz_io_p_1[378:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[17 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[17 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[17 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[12 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[12 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[12 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4[7 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[7 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[7 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[0 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[0 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[0 : 0];
  BADD_1125 NAFElements_adds_0 (
    .io_a   (NAFElements_adds_0_io_a[322:0]), //i
    .io_b   (NAFElements_adds_0_io_b[322:0]), //i
    .io_c   (1'b0                          ), //i
    .io_s   (NAFElements_adds_0_io_s[323:0]), //o
    .clk    (clk                           ), //i
    .resetn (resetn                        )  //i
  );
  BADD_1126 NAFElements_adds_1 (
    .io_a   (NAFElements_adds_1_io_a[332:0]), //i
    .io_b   (NAFElements_adds_1_io_b[332:0]), //i
    .io_c   (1'b0                          ), //i
    .io_s   (NAFElements_adds_1_io_s[333:0]), //o
    .clk    (clk                           ), //i
    .resetn (resetn                        )  //i
  );
  BADD_1127 NAFElements_adds_2 (
    .io_a   (NAFElements_adds_2_io_a[272:0]), //i
    .io_b   (NAFElements_adds_2_io_b[272:0]), //i
    .io_c   (1'b0                          ), //i
    .io_s   (NAFElements_adds_2_io_s[273:0]), //o
    .clk    (clk                           ), //i
    .resetn (resetn                        )  //i
  );
  BADD_1128 NAFElements_adds_3 (
    .io_a   (NAFElements_adds_3_io_a[189:0]), //i
    .io_b   (NAFElements_adds_3_io_b[189:0]), //i
    .io_c   (1'b1                          ), //i
    .io_s   (NAFElements_adds_3_io_s[190:0]), //o
    .clk    (clk                           ), //i
    .resetn (resetn                        )  //i
  );
  BADD_1129 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a[332:0]                                                                                                                                        ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[332:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[333:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1130 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_1[322:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[322:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[323:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1131 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[327:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[327:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[328:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1132 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_2[286:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[286:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[287:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1133 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_3[276:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[276:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[277:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1134 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[280:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[280:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[281:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1135 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[315:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[315:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[316:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_1136 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[253:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[253:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[254:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1137 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[234:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[234:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[235:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1138 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_4[239:0]                                                                                                                 ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[239:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[240:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1139 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[209:0]    ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1[209:0]), //i
    .io_c   (1'b0                                                                                                                                                       ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[210:0]    ), //o
    .clk    (clk                                                                                                                                                        ), //i
    .resetn (resetn                                                                                                                                                     )  //i
  );
  BADD_1140 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[170:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[170:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[171:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1141 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[176:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[176:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[177:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1142 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[214:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[214:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[215:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_1143 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[262:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[262:0]    ), //i
    .io_c   (1'b0                                                                                    ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[263:0]), //o
    .clk    (clk                                                                                     ), //i
    .resetn (resetn                                                                                  )  //i
  );
  BADD_1144 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_5[154:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[154:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[155:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1145 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[116:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[116:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[117:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_1146 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[136:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[136:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[137:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1147 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[106:0]    ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1[106:0]), //i
    .io_c   (1'b0                                                                                                                                                       ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[107:0]    ), //o
    .clk    (clk                                                                                                                                                        ), //i
    .resetn (resetn                                                                                                                                                     )  //i
  );
  BADD_1148 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[91:0]    ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1[91:0]), //i
    .io_c   (1'b0                                                                                                                                                      ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[92:0]    ), //o
    .clk    (clk                                                                                                                                                       ), //i
    .resetn (resetn                                                                                                                                                    )  //i
  );
  BADD_1149 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[101:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[101:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[102:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1150 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[111:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[111:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[112:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_1151 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[50:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[50:0]    ), //i
    .io_c   (1'b0                                                                                                                                                  ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[51:0]), //o
    .clk    (clk                                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                                )  //i
  );
  BADD_1152 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_6[42:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[42:0]    ), //i
    .io_c   (1'b0                                                                                                                                                  ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[43:0]), //o
    .clk    (clk                                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                                )  //i
  );
  BADD_1153 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_7[46:0]                                                                                                                 ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[46:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[47:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_1154 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[25:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[25:0]    ), //i
    .io_c   (1'b0                                                                                                                                                  ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[26:0]), //o
    .clk    (clk                                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                                )  //i
  );
  BADD_1155 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[15:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[15:0]    ), //i
    .io_c   (1'b0                                                                                                                                                  ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[16:0]), //o
    .clk    (clk                                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                                )  //i
  );
  BADD_1156 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[20:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[20:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[21:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_1157 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[31:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[31:0]    ), //i
    .io_c   (1'b0                                                                                                        ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[32:0]), //o
    .clk    (clk                                                                                                         ), //i
    .resetn (resetn                                                                                                      )  //i
  );
  BADD_1158 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[79:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[79:0]    ), //i
    .io_c   (1'b0                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[80:0]), //o
    .clk    (clk                                                                                    ), //i
    .resetn (resetn                                                                                 )  //i
  );
  BADD_1159 adder_posMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_a[162:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p[162:0]    ), //i
    .io_c   (1'b0                                                               ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_s[163:0]), //o
    .clk    (clk                                                                ), //i
    .resetn (resetn                                                             )  //i
  );
  BADD_1160 adder_posMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_add_add_io_a[4:0]    ), //i
    .io_b   (adder_posMUL_multiElements_msbMUL_p_delay_5[4:0]), //i
    .io_c   (1'b0                                            ), //i
    .io_s   (adder_posMUL_multiElements_add_add_io_s[5:0]    ), //o
    .clk    (clk                                             ), //i
    .resetn (resetn                                          )  //i
  );
  BADD_1161 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[267:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[267:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[268:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1162 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[225:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[225:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[226:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1163 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[258:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[258:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[259:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_1164 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_8[205:0]                                                                                                                 ), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[205:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[206:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1165 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[194:0]    ), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1[194:0]), //i
    .io_c   (1'b0                                                                                                                                  ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[195:0]    ), //o
    .clk    (clk                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                )  //i
  );
  BADD_1166 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[200:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[200:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[201:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_1167 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[220:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[220:0]    ), //i
    .io_c   (1'b0                                                                                    ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[221:0]), //o
    .clk    (clk                                                                                     ), //i
    .resetn (resetn                                                                                  )  //i
  );
  BADD_1168 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[182:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[182:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[183:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1169 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[150:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[150:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[151:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1170 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[166:0]    ), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1[166:0]), //i
    .io_c   (1'b0                                                                                                             ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[167:0]    ), //o
    .clk    (clk                                                                                                              ), //i
    .resetn (resetn                                                                                                           )  //i
  );
  BADD_1171 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[141:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[141:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[142:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1172 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[125:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[125:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[126:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_1173 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[129:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[129:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[130:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_1174 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[145:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[145:0]    ), //i
    .io_c   (1'b0                                                                                    ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[146:0]), //o
    .clk    (clk                                                                                     ), //i
    .resetn (resetn                                                                                  )  //i
  );
  BADD_1175 adder_negMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_a[189:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p[189:0]    ), //i
    .io_c   (1'b0                                                               ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_s[190:0]), //o
    .clk    (clk                                                                ), //i
    .resetn (resetn                                                             )  //i
  );
  BADD_1176 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_9[96:0]                                                                                                                 ), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[96:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[97:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_1177 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[74:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[74:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[75:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_1178 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[84:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[84:0]    ), //i
    .io_c   (1'b0                                                                                                        ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[85:0]), //o
    .clk    (clk                                                                                                         ), //i
    .resetn (resetn                                                                                                      )  //i
  );
  BADD_1179 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[63:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[64:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_1180 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[54:0]    ), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1[54:0]), //i
    .io_c   (1'b0                                                                                                                                 ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[55:0]    ), //o
    .clk    (clk                                                                                                                                  ), //i
    .resetn (resetn                                                                                                                               )  //i
  );
  BADD_1181 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[58:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[58:0]    ), //i
    .io_c   (1'b0                                                                                                        ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[59:0]), //o
    .clk    (clk                                                                                                         ), //i
    .resetn (resetn                                                                                                      )  //i
  );
  BADD_1182 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[68:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[68:0]    ), //i
    .io_c   (1'b0                                                                                   ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[69:0]), //o
    .clk    (clk                                                                                    ), //i
    .resetn (resetn                                                                                 )  //i
  );
  BADD_1183 adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_10[9:0]                                                                       ), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[9:0]     ), //i
    .io_c   (1'b0                                                                                   ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[10:0]), //o
    .clk    (clk                                                                                    ), //i
    .resetn (resetn                                                                                 )  //i
  );
  BADD_1184 adder_negMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_a[36:0]    ), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_2[36:0]), //i
    .io_c   (1'b0                                                                  ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_s[37:0]    ), //o
    .clk    (clk                                                                   ), //i
    .resetn (resetn                                                                )  //i
  );
  BADD_1185 adder_negMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_add_add_io_a[120:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_p[120:0]    ), //i
    .io_c   (1'b0                                          ), //i
    .io_s   (adder_negMUL_multiElements_add_add_io_s[121:0]), //o
    .clk    (clk                                           ), //i
    .resetn (resetn                                        )  //i
  );
  BADD_1186 adder_add (
    .io_a   (adder_posMUL_p[378:0]), //i
    .io_b   (adder_add_io_b[378:0]), //i
    .io_c   (1'b1                 ), //i
    .io_s   (adder_add_io_s[379:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign NAFElements_adds_0_io_a = _zz_io_a_11[322:0];
  assign NAFElements_adds_0_io_b = io_a[322:0];
  assign NAFElements_adds_1_io_a = _zz_io_a_12[332:0];
  assign NAFElements_adds_1_io_b = io_a[332:0];
  assign NAFElements_adds_2_io_a = _zz_io_a_13[272:0];
  assign NAFElements_adds_2_io_b = io_a[272:0];
  assign NAFElements_adds_3_io_a = _zz_io_a_14[189:0];
  assign NAFElements_adds_3_io_b = io_a[189:0];
  assign _zz_NAFElements_sums_0 = {1'd0, io_a};
  assign NAFElements_sums_0 = {_zz_NAFElements_sums_0_15,{_zz_NAFElements_sums_0_10,{_zz_NAFElements_sums_0_6,{_zz_NAFElements_sums_0_3,{_zz_NAFElements_sums_0_1,_zz_NAFElements_sums_0[63 : 0]}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_adds_0_io_s[322:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_adds_1_io_s[332:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_adds_2_io_s[272:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_adds_3_io_s[189:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 320],{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[319 : 256],{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[255 : 192],{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128],{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64],_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0]}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[255 : 192];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[319 : 256];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[332 : 320],{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6[17 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5[17 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14}}}}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[45 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 46] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[332:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[327:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[255 : 192];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[319 : 256];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[327 : 320],{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5[12 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[12 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13}}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[255 : 192];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[319 : 256];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[322 : 320],{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6[7 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5[7 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14}}}}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[327 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[322:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 51);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[50 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 51] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[327:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[315:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[255 : 192];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[315 : 256];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5[0 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[0 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[286:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[255 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7}}}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[28 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[315 : 29] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[286:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[280:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[255 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[276:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[255 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7}}}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[3 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[280 : 4] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[276:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 35);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[34 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[315 : 35] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[280:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 63);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[62 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 63] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[315:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[262:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[255 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_sums_0[253:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[253 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7}}}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 9);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[8 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[262 : 9] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[253:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[239:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[234:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8}}}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[239 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[234:0];
  end

  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[22 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[262 : 23] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[239:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[214:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_sums_0[209:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8}}}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[214 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[209:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[176:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[170:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9}}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 6);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[5 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[176 : 6] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[170:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 38);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[37 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[214 : 38] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[176:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 48);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[47 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[262 : 48] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[214:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 116);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[115 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 116] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[262:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[162:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[154:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[7 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[162 : 8] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[154:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[136:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[116:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 20);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[19 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[136 : 20] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[116:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 26);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[25 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[162 : 26] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[136:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[111:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_sums_0[106:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[111 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[106:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[101:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_sums_0[91:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 10);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[9 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[101 : 10] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[91:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 10);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[9 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[111 : 10] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[101:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 51);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[50 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[162 : 51] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[111:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[79:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 29);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[28 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[79 : 29] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[50:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[3 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[46 : 4] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[42:0];
  end

  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[32 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[79 : 33] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[46:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 6);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[5 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[31 : 6] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[25:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[20 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[15:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 11);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[10 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[31 : 11] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[20:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 48);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[47 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[79 : 48] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[31:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 83);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p[82 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p[162 : 83] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[79:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 216);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_p[215 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_p[378 : 216] = adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_s[162:0];
  end

  assign adder_posMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_msbMUL_p_4;
  assign adder_posMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_p >>> 374);
  always @(*) begin
    adder_posMUL_p[373 : 0] = _zz_adder_posMUL_p;
    adder_posMUL_p[378 : 374] = adder_posMUL_multiElements_add_add_io_s[4:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[191 : 128];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[255 : 192];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8}}}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[267:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[255 : 192];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7}}}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[272 : 5] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[267:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[258:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[255 : 192];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7}}}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[225:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8}}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 33);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[32 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[258 : 33] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[225:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 14);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[13 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[272 : 14] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[258:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[220:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8}}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[205:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8}}}};
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[14 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[220 : 15] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[205:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[200:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8}}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_sums_0[194:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8}}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 6);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[5 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[200 : 6] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[194:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 20);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[19 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[220 : 20] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[200:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 52);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[51 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[272 : 52] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[220:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[189 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[182:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 7);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[6 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[189 : 7] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[182:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[166:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_sums_0[150:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 16);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[15 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[166 : 16] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[150:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 23);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[22 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[189 : 23] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[166:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[145:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[141:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 4);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[145 : 4] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[141:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[129:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[125:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[125 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 4);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[3 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[129 : 4] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[125:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 16);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[15 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[145 : 16] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[129:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 44);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p[43 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p[189 : 44] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[145:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 83);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_p[82 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_p[272 : 83] = adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_s[189:0];
  end

  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[120:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[96:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10}};
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[23 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[120 : 24] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[96:0];
  end

  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[84:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[74:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10}};
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 10);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[9 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[84 : 10] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[74:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 36);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[35 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[120 : 36] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[84:0];
  end

  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[68:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9};
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[68 : 5] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[63:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 4);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[3 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[58 : 4] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[54:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 10);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[9 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[68 : 10] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[58:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 52);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p[51 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p[120 : 52] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[68:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  assign adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p[26 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p[36 : 27] = adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[9:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 84);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_p[83 : 0] = _zz_adder_negMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_p[120 : 84] = adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_s[36:0];
  end

  assign adder_negMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_p >>> 152);
  always @(*) begin
    adder_negMUL_p[151 : 0] = _zz_adder_negMUL_p;
    adder_negMUL_p[272 : 152] = adder_negMUL_multiElements_add_add_io_s[120:0];
  end

  assign adder_add_io_b = ({106'd0,adder_negMUL_p_delay_1} <<< 106);
  assign io_p[378 : 0] = _zz_io_p;
  always @(posedge clk) begin
    _zz_NAFElements_sums_0_1 <= _zz_NAFElements_sums_0[127 : 64];
    _zz_NAFElements_sums_0_2 <= _zz_NAFElements_sums_0[191 : 128];
    _zz_NAFElements_sums_0_3 <= _zz_NAFElements_sums_0_2;
    _zz_NAFElements_sums_0_4 <= _zz_NAFElements_sums_0[255 : 192];
    _zz_NAFElements_sums_0_5 <= _zz_NAFElements_sums_0_4;
    _zz_NAFElements_sums_0_6 <= _zz_NAFElements_sums_0_5;
    _zz_NAFElements_sums_0_7 <= _zz_NAFElements_sums_0[319 : 256];
    _zz_NAFElements_sums_0_8 <= _zz_NAFElements_sums_0_7;
    _zz_NAFElements_sums_0_9 <= _zz_NAFElements_sums_0_8;
    _zz_NAFElements_sums_0_10 <= _zz_NAFElements_sums_0_9;
    _zz_NAFElements_sums_0_11 <= _zz_NAFElements_sums_0[378 : 320];
    _zz_NAFElements_sums_0_12 <= _zz_NAFElements_sums_0_11;
    _zz_NAFElements_sums_0_13 <= _zz_NAFElements_sums_0_12;
    _zz_NAFElements_sums_0_14 <= _zz_NAFElements_sums_0_13;
    _zz_NAFElements_sums_0_15 <= _zz_NAFElements_sums_0_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 18];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 18];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[63 : 18];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5[63 : 18];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6[63 : 18];
    _zz_io_a <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 46);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[45 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 8];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 8];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4[63 : 8];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5[63 : 8];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6[63 : 8];
    _zz_io_a_1 <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 5);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[50 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[63 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5[59 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 36];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[35 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 36];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[35 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 36];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[35 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[63 : 36];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[35 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[286 : 256];
    _zz_io_a_2 <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 29);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[28 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 30];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[29 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 30];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[29 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 30];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[29 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[63 : 30];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[29 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[280 : 256];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 26];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 26];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 26];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4[63 : 26];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[276 : 256];
    _zz_io_a_3 <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 4);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[34 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[62 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 12];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[11 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 12];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[11 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 12];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[11 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[63 : 12];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[11 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[262 : 256];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 3];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[2 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 3];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[2 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 3];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[2 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[61 : 3];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[2 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[8 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 53];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[52 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 53];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[52 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 53];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[52 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[239 : 192];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[234 : 192];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_io_a_4 <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 23);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[22 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 28];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[27 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 28];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[27 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 28];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[27 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[214 : 192];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 23];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[22 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 23];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[22 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 23];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[22 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[209 : 192];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1 <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 54];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[53 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 54];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[53 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[176 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[170 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[5 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[37 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[115 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 40];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[39 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 40];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[39 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[162 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 32];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[31 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 32];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[31 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[154 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
    _zz_io_a_5 <= (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 8);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[7 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 14];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[13 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 14];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[13 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[136 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 58];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[57 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[116 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[19 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 53];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[52 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[111 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[106 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1 <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 43];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[42 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[101 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 33];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[32 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[91 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1 <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[9 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[9 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[50 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 21];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[20 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[79 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[50 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[28 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[46 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[42 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_io_a_6 <= (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 4);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_io_a_7 <= (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 33);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[32 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[31 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[5 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[20 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[15 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[10 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[82 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[215 : 0];
    _zz_adder_posMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_msbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_msbMUL_p_3;
    adder_posMUL_multiElements_msbMUL_p_delay_1 <= adder_posMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_msbMUL_p_delay_2 <= adder_posMUL_multiElements_msbMUL_p_delay_1;
    adder_posMUL_multiElements_msbMUL_p_delay_3 <= adder_posMUL_multiElements_msbMUL_p_delay_2;
    adder_posMUL_multiElements_msbMUL_p_delay_4 <= adder_posMUL_multiElements_msbMUL_p_delay_3;
    adder_posMUL_multiElements_msbMUL_p_delay_5 <= adder_posMUL_multiElements_msbMUL_p_delay_4;
    _zz_adder_posMUL_p <= adder_posMUL_multiElements_lsbMUL_p[373 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 22];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[21 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 22];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[21 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[63 : 22];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[21 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5[63 : 22];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5[21 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[272 : 256];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 17];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[16 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 17];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[16 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 17];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[16 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[63 : 17];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[16 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[267 : 256];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[258 : 256];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 39];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[38 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 39];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[38 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 39];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[38 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[225 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[32 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[13 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 34];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[33 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 34];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[33 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 34];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[33 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[220 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[205 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
    _zz_io_a_8 <= (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 15);
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[14 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 14];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[13 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 14];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[13 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 14];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[13 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[200 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[194 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1 <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[5 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[19 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[51 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[61 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 60];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[59 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 60];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[59 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[182 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[6 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 44];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[43 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 44];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[43 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[166 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 28];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[27 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 28];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[27 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[150 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[15 : 0];
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1 <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[22 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 23];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[22 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 23];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[22 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[145 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[141 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 7];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[6 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 7];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[6 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[129 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[61 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[15 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[43 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[82 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 62];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[61 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[120 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 38];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[37 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[96 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
    _zz_io_a_9 <= (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 24);
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[23 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 26];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[25 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[84 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 16];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[15 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[74 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[9 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[35 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 10];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[9 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[68 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 5];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[4 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[58 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[54 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1 <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[9 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[51 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[36 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[9 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_io_a_10 <= (adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 27);
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[26 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1 <= adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_2 <= adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
    _zz_adder_negMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p[83 : 0];
    _zz_adder_negMUL_p <= adder_negMUL_multiElements_lsbMUL_p[151 : 0];
    adder_negMUL_p_delay_1 <= adder_negMUL_p;
  end


endmodule

module KaratsubaMUL_35 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  output     [755:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [47:0]   core_io_a_0;
  wire       [47:0]   core_io_a_1;
  wire       [47:0]   core_io_a_2;
  wire       [47:0]   core_io_a_3;
  wire       [47:0]   core_io_a_4;
  wire       [47:0]   core_io_a_5;
  wire       [47:0]   core_io_a_6;
  wire       [47:0]   core_io_a_7;
  wire       [47:0]   core_io_b_0;
  wire       [47:0]   core_io_b_1;
  wire       [47:0]   core_io_b_2;
  wire       [47:0]   core_io_b_3;
  wire       [47:0]   core_io_b_4;
  wire       [47:0]   core_io_b_5;
  wire       [47:0]   core_io_b_6;
  wire       [47:0]   core_io_b_7;
  wire       [767:0]  core_io_p;
  wire       [47:0]   _zz_io_p_121;
  wire       [239:0]  _zz_io_p_122;
  wire       [383:0]  a;
  wire       [383:0]  b;
  wire       [335:0]  _zz_io_a_0;
  wire       [335:0]  _zz_io_b_0;
  wire       [755:0]  _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;
  reg        [47:0]   _zz_io_p_4;
  reg        [47:0]   _zz_io_p_5;
  reg        [47:0]   _zz_io_p_6;
  reg        [47:0]   _zz_io_p_7;
  reg        [47:0]   _zz_io_p_8;
  reg        [47:0]   _zz_io_p_9;
  reg        [47:0]   _zz_io_p_10;
  reg        [47:0]   _zz_io_p_11;
  reg        [47:0]   _zz_io_p_12;
  reg        [47:0]   _zz_io_p_13;
  reg        [47:0]   _zz_io_p_14;
  reg        [47:0]   _zz_io_p_15;
  reg        [47:0]   _zz_io_p_16;
  reg        [47:0]   _zz_io_p_17;
  reg        [47:0]   _zz_io_p_18;
  reg        [47:0]   _zz_io_p_19;
  reg        [47:0]   _zz_io_p_20;
  reg        [47:0]   _zz_io_p_21;
  reg        [47:0]   _zz_io_p_22;
  reg        [47:0]   _zz_io_p_23;
  reg        [47:0]   _zz_io_p_24;
  reg        [47:0]   _zz_io_p_25;
  reg        [47:0]   _zz_io_p_26;
  reg        [47:0]   _zz_io_p_27;
  reg        [47:0]   _zz_io_p_28;
  reg        [47:0]   _zz_io_p_29;
  reg        [47:0]   _zz_io_p_30;
  reg        [47:0]   _zz_io_p_31;
  reg        [47:0]   _zz_io_p_32;
  reg        [47:0]   _zz_io_p_33;
  reg        [47:0]   _zz_io_p_34;
  reg        [47:0]   _zz_io_p_35;
  reg        [47:0]   _zz_io_p_36;
  reg        [47:0]   _zz_io_p_37;
  reg        [47:0]   _zz_io_p_38;
  reg        [47:0]   _zz_io_p_39;
  reg        [47:0]   _zz_io_p_40;
  reg        [47:0]   _zz_io_p_41;
  reg        [47:0]   _zz_io_p_42;
  reg        [47:0]   _zz_io_p_43;
  reg        [47:0]   _zz_io_p_44;
  reg        [47:0]   _zz_io_p_45;
  reg        [47:0]   _zz_io_p_46;
  reg        [47:0]   _zz_io_p_47;
  reg        [47:0]   _zz_io_p_48;
  reg        [47:0]   _zz_io_p_49;
  reg        [47:0]   _zz_io_p_50;
  reg        [47:0]   _zz_io_p_51;
  reg        [47:0]   _zz_io_p_52;
  reg        [47:0]   _zz_io_p_53;
  reg        [47:0]   _zz_io_p_54;
  reg        [47:0]   _zz_io_p_55;
  reg        [47:0]   _zz_io_p_56;
  reg        [47:0]   _zz_io_p_57;
  reg        [47:0]   _zz_io_p_58;
  reg        [47:0]   _zz_io_p_59;
  reg        [47:0]   _zz_io_p_60;
  reg        [47:0]   _zz_io_p_61;
  reg        [47:0]   _zz_io_p_62;
  reg        [47:0]   _zz_io_p_63;
  reg        [47:0]   _zz_io_p_64;
  reg        [47:0]   _zz_io_p_65;
  reg        [47:0]   _zz_io_p_66;
  reg        [47:0]   _zz_io_p_67;
  reg        [47:0]   _zz_io_p_68;
  reg        [47:0]   _zz_io_p_69;
  reg        [47:0]   _zz_io_p_70;
  reg        [47:0]   _zz_io_p_71;
  reg        [47:0]   _zz_io_p_72;
  reg        [47:0]   _zz_io_p_73;
  reg        [47:0]   _zz_io_p_74;
  reg        [47:0]   _zz_io_p_75;
  reg        [47:0]   _zz_io_p_76;
  reg        [47:0]   _zz_io_p_77;
  reg        [47:0]   _zz_io_p_78;
  reg        [47:0]   _zz_io_p_79;
  reg        [47:0]   _zz_io_p_80;
  reg        [47:0]   _zz_io_p_81;
  reg        [47:0]   _zz_io_p_82;
  reg        [47:0]   _zz_io_p_83;
  reg        [47:0]   _zz_io_p_84;
  reg        [47:0]   _zz_io_p_85;
  reg        [47:0]   _zz_io_p_86;
  reg        [47:0]   _zz_io_p_87;
  reg        [47:0]   _zz_io_p_88;
  reg        [47:0]   _zz_io_p_89;
  reg        [47:0]   _zz_io_p_90;
  reg        [47:0]   _zz_io_p_91;
  reg        [47:0]   _zz_io_p_92;
  reg        [47:0]   _zz_io_p_93;
  reg        [47:0]   _zz_io_p_94;
  reg        [47:0]   _zz_io_p_95;
  reg        [47:0]   _zz_io_p_96;
  reg        [47:0]   _zz_io_p_97;
  reg        [47:0]   _zz_io_p_98;
  reg        [47:0]   _zz_io_p_99;
  reg        [47:0]   _zz_io_p_100;
  reg        [47:0]   _zz_io_p_101;
  reg        [47:0]   _zz_io_p_102;
  reg        [47:0]   _zz_io_p_103;
  reg        [47:0]   _zz_io_p_104;
  reg        [47:0]   _zz_io_p_105;
  reg        [47:0]   _zz_io_p_106;
  reg        [47:0]   _zz_io_p_107;
  reg        [47:0]   _zz_io_p_108;
  reg        [47:0]   _zz_io_p_109;
  reg        [47:0]   _zz_io_p_110;
  reg        [47:0]   _zz_io_p_111;
  reg        [47:0]   _zz_io_p_112;
  reg        [47:0]   _zz_io_p_113;
  reg        [47:0]   _zz_io_p_114;
  reg        [47:0]   _zz_io_p_115;
  reg        [47:0]   _zz_io_p_116;
  reg        [47:0]   _zz_io_p_117;
  reg        [47:0]   _zz_io_p_118;
  reg        [47:0]   _zz_io_p_119;
  reg        [47:0]   _zz_io_p_120;

  assign _zz_io_p_121 = _zz_io_p_75;
  assign _zz_io_p_122 = {_zz_io_p_65,{_zz_io_p_54,{_zz_io_p_42,{_zz_io_p_29,_zz_io_p_15}}}};
  KaratsubaCore_35 core (
    .io_a_0 (core_io_a_0[47:0]), //i
    .io_a_1 (core_io_a_1[47:0]), //i
    .io_a_2 (core_io_a_2[47:0]), //i
    .io_a_3 (core_io_a_3[47:0]), //i
    .io_a_4 (core_io_a_4[47:0]), //i
    .io_a_5 (core_io_a_5[47:0]), //i
    .io_a_6 (core_io_a_6[47:0]), //i
    .io_a_7 (core_io_a_7[47:0]), //i
    .io_b_0 (core_io_b_0[47:0]), //i
    .io_b_1 (core_io_b_1[47:0]), //i
    .io_b_2 (core_io_b_2[47:0]), //i
    .io_b_3 (core_io_b_3[47:0]), //i
    .io_b_4 (core_io_b_4[47:0]), //i
    .io_b_5 (core_io_b_5[47:0]), //i
    .io_b_6 (core_io_b_6[47:0]), //i
    .io_b_7 (core_io_b_7[47:0]), //i
    .io_p   (core_io_p[767:0] ), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  assign a = {6'd0, io_a};
  assign b = {6'd0, io_b};
  assign _zz_io_a_0 = a[335:0];
  assign core_io_a_0 = _zz_io_a_0[47 : 0];
  assign core_io_a_1 = _zz_io_a_0[95 : 48];
  assign core_io_a_2 = _zz_io_a_0[143 : 96];
  assign core_io_a_3 = _zz_io_a_0[191 : 144];
  assign core_io_a_4 = _zz_io_a_0[239 : 192];
  assign core_io_a_5 = _zz_io_a_0[287 : 240];
  assign core_io_a_6 = _zz_io_a_0[335 : 288];
  assign core_io_a_7 = (a >>> 336);
  assign _zz_io_b_0 = b[335:0];
  assign core_io_b_0 = _zz_io_b_0[47 : 0];
  assign core_io_b_1 = _zz_io_b_0[95 : 48];
  assign core_io_b_2 = _zz_io_b_0[143 : 96];
  assign core_io_b_3 = _zz_io_b_0[191 : 144];
  assign core_io_b_4 = _zz_io_b_0[239 : 192];
  assign core_io_b_5 = _zz_io_b_0[287 : 240];
  assign core_io_b_6 = _zz_io_b_0[335 : 288];
  assign core_io_b_7 = (b >>> 336);
  assign _zz_io_p = core_io_p[755:0];
  assign io_p = {_zz_io_p[755 : 720],{_zz_io_p_120,{_zz_io_p_119,{_zz_io_p_117,{_zz_io_p_114,{_zz_io_p_110,{_zz_io_p_105,{_zz_io_p_99,{_zz_io_p_92,{_zz_io_p_84,{_zz_io_p_121,_zz_io_p_122}}}}}}}}}}};
  always @(posedge clk) begin
    _zz_io_p_1 <= _zz_io_p[47 : 0];
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= _zz_io_p_2;
    _zz_io_p_4 <= _zz_io_p_3;
    _zz_io_p_5 <= _zz_io_p_4;
    _zz_io_p_6 <= _zz_io_p_5;
    _zz_io_p_7 <= _zz_io_p_6;
    _zz_io_p_8 <= _zz_io_p_7;
    _zz_io_p_9 <= _zz_io_p_8;
    _zz_io_p_10 <= _zz_io_p_9;
    _zz_io_p_11 <= _zz_io_p_10;
    _zz_io_p_12 <= _zz_io_p_11;
    _zz_io_p_13 <= _zz_io_p_12;
    _zz_io_p_14 <= _zz_io_p_13;
    _zz_io_p_15 <= _zz_io_p_14;
    _zz_io_p_16 <= _zz_io_p[95 : 48];
    _zz_io_p_17 <= _zz_io_p_16;
    _zz_io_p_18 <= _zz_io_p_17;
    _zz_io_p_19 <= _zz_io_p_18;
    _zz_io_p_20 <= _zz_io_p_19;
    _zz_io_p_21 <= _zz_io_p_20;
    _zz_io_p_22 <= _zz_io_p_21;
    _zz_io_p_23 <= _zz_io_p_22;
    _zz_io_p_24 <= _zz_io_p_23;
    _zz_io_p_25 <= _zz_io_p_24;
    _zz_io_p_26 <= _zz_io_p_25;
    _zz_io_p_27 <= _zz_io_p_26;
    _zz_io_p_28 <= _zz_io_p_27;
    _zz_io_p_29 <= _zz_io_p_28;
    _zz_io_p_30 <= _zz_io_p[143 : 96];
    _zz_io_p_31 <= _zz_io_p_30;
    _zz_io_p_32 <= _zz_io_p_31;
    _zz_io_p_33 <= _zz_io_p_32;
    _zz_io_p_34 <= _zz_io_p_33;
    _zz_io_p_35 <= _zz_io_p_34;
    _zz_io_p_36 <= _zz_io_p_35;
    _zz_io_p_37 <= _zz_io_p_36;
    _zz_io_p_38 <= _zz_io_p_37;
    _zz_io_p_39 <= _zz_io_p_38;
    _zz_io_p_40 <= _zz_io_p_39;
    _zz_io_p_41 <= _zz_io_p_40;
    _zz_io_p_42 <= _zz_io_p_41;
    _zz_io_p_43 <= _zz_io_p[191 : 144];
    _zz_io_p_44 <= _zz_io_p_43;
    _zz_io_p_45 <= _zz_io_p_44;
    _zz_io_p_46 <= _zz_io_p_45;
    _zz_io_p_47 <= _zz_io_p_46;
    _zz_io_p_48 <= _zz_io_p_47;
    _zz_io_p_49 <= _zz_io_p_48;
    _zz_io_p_50 <= _zz_io_p_49;
    _zz_io_p_51 <= _zz_io_p_50;
    _zz_io_p_52 <= _zz_io_p_51;
    _zz_io_p_53 <= _zz_io_p_52;
    _zz_io_p_54 <= _zz_io_p_53;
    _zz_io_p_55 <= _zz_io_p[239 : 192];
    _zz_io_p_56 <= _zz_io_p_55;
    _zz_io_p_57 <= _zz_io_p_56;
    _zz_io_p_58 <= _zz_io_p_57;
    _zz_io_p_59 <= _zz_io_p_58;
    _zz_io_p_60 <= _zz_io_p_59;
    _zz_io_p_61 <= _zz_io_p_60;
    _zz_io_p_62 <= _zz_io_p_61;
    _zz_io_p_63 <= _zz_io_p_62;
    _zz_io_p_64 <= _zz_io_p_63;
    _zz_io_p_65 <= _zz_io_p_64;
    _zz_io_p_66 <= _zz_io_p[287 : 240];
    _zz_io_p_67 <= _zz_io_p_66;
    _zz_io_p_68 <= _zz_io_p_67;
    _zz_io_p_69 <= _zz_io_p_68;
    _zz_io_p_70 <= _zz_io_p_69;
    _zz_io_p_71 <= _zz_io_p_70;
    _zz_io_p_72 <= _zz_io_p_71;
    _zz_io_p_73 <= _zz_io_p_72;
    _zz_io_p_74 <= _zz_io_p_73;
    _zz_io_p_75 <= _zz_io_p_74;
    _zz_io_p_76 <= _zz_io_p[335 : 288];
    _zz_io_p_77 <= _zz_io_p_76;
    _zz_io_p_78 <= _zz_io_p_77;
    _zz_io_p_79 <= _zz_io_p_78;
    _zz_io_p_80 <= _zz_io_p_79;
    _zz_io_p_81 <= _zz_io_p_80;
    _zz_io_p_82 <= _zz_io_p_81;
    _zz_io_p_83 <= _zz_io_p_82;
    _zz_io_p_84 <= _zz_io_p_83;
    _zz_io_p_85 <= _zz_io_p[383 : 336];
    _zz_io_p_86 <= _zz_io_p_85;
    _zz_io_p_87 <= _zz_io_p_86;
    _zz_io_p_88 <= _zz_io_p_87;
    _zz_io_p_89 <= _zz_io_p_88;
    _zz_io_p_90 <= _zz_io_p_89;
    _zz_io_p_91 <= _zz_io_p_90;
    _zz_io_p_92 <= _zz_io_p_91;
    _zz_io_p_93 <= _zz_io_p[431 : 384];
    _zz_io_p_94 <= _zz_io_p_93;
    _zz_io_p_95 <= _zz_io_p_94;
    _zz_io_p_96 <= _zz_io_p_95;
    _zz_io_p_97 <= _zz_io_p_96;
    _zz_io_p_98 <= _zz_io_p_97;
    _zz_io_p_99 <= _zz_io_p_98;
    _zz_io_p_100 <= _zz_io_p[479 : 432];
    _zz_io_p_101 <= _zz_io_p_100;
    _zz_io_p_102 <= _zz_io_p_101;
    _zz_io_p_103 <= _zz_io_p_102;
    _zz_io_p_104 <= _zz_io_p_103;
    _zz_io_p_105 <= _zz_io_p_104;
    _zz_io_p_106 <= _zz_io_p[527 : 480];
    _zz_io_p_107 <= _zz_io_p_106;
    _zz_io_p_108 <= _zz_io_p_107;
    _zz_io_p_109 <= _zz_io_p_108;
    _zz_io_p_110 <= _zz_io_p_109;
    _zz_io_p_111 <= _zz_io_p[575 : 528];
    _zz_io_p_112 <= _zz_io_p_111;
    _zz_io_p_113 <= _zz_io_p_112;
    _zz_io_p_114 <= _zz_io_p_113;
    _zz_io_p_115 <= _zz_io_p[623 : 576];
    _zz_io_p_116 <= _zz_io_p_115;
    _zz_io_p_117 <= _zz_io_p_116;
    _zz_io_p_118 <= _zz_io_p[671 : 624];
    _zz_io_p_119 <= _zz_io_p_118;
    _zz_io_p_120 <= _zz_io_p[719 : 672];
  end


endmodule

module KaratsubaMUL_34 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  output     [753:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [47:0]   core_io_a_0;
  wire       [47:0]   core_io_a_1;
  wire       [47:0]   core_io_a_2;
  wire       [47:0]   core_io_a_3;
  wire       [47:0]   core_io_a_4;
  wire       [47:0]   core_io_a_5;
  wire       [47:0]   core_io_a_6;
  wire       [47:0]   core_io_a_7;
  wire       [47:0]   core_io_b_0;
  wire       [47:0]   core_io_b_1;
  wire       [47:0]   core_io_b_2;
  wire       [47:0]   core_io_b_3;
  wire       [47:0]   core_io_b_4;
  wire       [47:0]   core_io_b_5;
  wire       [47:0]   core_io_b_6;
  wire       [47:0]   core_io_b_7;
  wire       [767:0]  core_io_p;
  wire       [47:0]   _zz_io_p_121;
  wire       [239:0]  _zz_io_p_122;
  wire       [383:0]  a;
  wire       [383:0]  b;
  wire       [335:0]  _zz_io_a_0;
  wire       [335:0]  _zz_io_b_0;
  wire       [753:0]  _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;
  reg        [47:0]   _zz_io_p_4;
  reg        [47:0]   _zz_io_p_5;
  reg        [47:0]   _zz_io_p_6;
  reg        [47:0]   _zz_io_p_7;
  reg        [47:0]   _zz_io_p_8;
  reg        [47:0]   _zz_io_p_9;
  reg        [47:0]   _zz_io_p_10;
  reg        [47:0]   _zz_io_p_11;
  reg        [47:0]   _zz_io_p_12;
  reg        [47:0]   _zz_io_p_13;
  reg        [47:0]   _zz_io_p_14;
  reg        [47:0]   _zz_io_p_15;
  reg        [47:0]   _zz_io_p_16;
  reg        [47:0]   _zz_io_p_17;
  reg        [47:0]   _zz_io_p_18;
  reg        [47:0]   _zz_io_p_19;
  reg        [47:0]   _zz_io_p_20;
  reg        [47:0]   _zz_io_p_21;
  reg        [47:0]   _zz_io_p_22;
  reg        [47:0]   _zz_io_p_23;
  reg        [47:0]   _zz_io_p_24;
  reg        [47:0]   _zz_io_p_25;
  reg        [47:0]   _zz_io_p_26;
  reg        [47:0]   _zz_io_p_27;
  reg        [47:0]   _zz_io_p_28;
  reg        [47:0]   _zz_io_p_29;
  reg        [47:0]   _zz_io_p_30;
  reg        [47:0]   _zz_io_p_31;
  reg        [47:0]   _zz_io_p_32;
  reg        [47:0]   _zz_io_p_33;
  reg        [47:0]   _zz_io_p_34;
  reg        [47:0]   _zz_io_p_35;
  reg        [47:0]   _zz_io_p_36;
  reg        [47:0]   _zz_io_p_37;
  reg        [47:0]   _zz_io_p_38;
  reg        [47:0]   _zz_io_p_39;
  reg        [47:0]   _zz_io_p_40;
  reg        [47:0]   _zz_io_p_41;
  reg        [47:0]   _zz_io_p_42;
  reg        [47:0]   _zz_io_p_43;
  reg        [47:0]   _zz_io_p_44;
  reg        [47:0]   _zz_io_p_45;
  reg        [47:0]   _zz_io_p_46;
  reg        [47:0]   _zz_io_p_47;
  reg        [47:0]   _zz_io_p_48;
  reg        [47:0]   _zz_io_p_49;
  reg        [47:0]   _zz_io_p_50;
  reg        [47:0]   _zz_io_p_51;
  reg        [47:0]   _zz_io_p_52;
  reg        [47:0]   _zz_io_p_53;
  reg        [47:0]   _zz_io_p_54;
  reg        [47:0]   _zz_io_p_55;
  reg        [47:0]   _zz_io_p_56;
  reg        [47:0]   _zz_io_p_57;
  reg        [47:0]   _zz_io_p_58;
  reg        [47:0]   _zz_io_p_59;
  reg        [47:0]   _zz_io_p_60;
  reg        [47:0]   _zz_io_p_61;
  reg        [47:0]   _zz_io_p_62;
  reg        [47:0]   _zz_io_p_63;
  reg        [47:0]   _zz_io_p_64;
  reg        [47:0]   _zz_io_p_65;
  reg        [47:0]   _zz_io_p_66;
  reg        [47:0]   _zz_io_p_67;
  reg        [47:0]   _zz_io_p_68;
  reg        [47:0]   _zz_io_p_69;
  reg        [47:0]   _zz_io_p_70;
  reg        [47:0]   _zz_io_p_71;
  reg        [47:0]   _zz_io_p_72;
  reg        [47:0]   _zz_io_p_73;
  reg        [47:0]   _zz_io_p_74;
  reg        [47:0]   _zz_io_p_75;
  reg        [47:0]   _zz_io_p_76;
  reg        [47:0]   _zz_io_p_77;
  reg        [47:0]   _zz_io_p_78;
  reg        [47:0]   _zz_io_p_79;
  reg        [47:0]   _zz_io_p_80;
  reg        [47:0]   _zz_io_p_81;
  reg        [47:0]   _zz_io_p_82;
  reg        [47:0]   _zz_io_p_83;
  reg        [47:0]   _zz_io_p_84;
  reg        [47:0]   _zz_io_p_85;
  reg        [47:0]   _zz_io_p_86;
  reg        [47:0]   _zz_io_p_87;
  reg        [47:0]   _zz_io_p_88;
  reg        [47:0]   _zz_io_p_89;
  reg        [47:0]   _zz_io_p_90;
  reg        [47:0]   _zz_io_p_91;
  reg        [47:0]   _zz_io_p_92;
  reg        [47:0]   _zz_io_p_93;
  reg        [47:0]   _zz_io_p_94;
  reg        [47:0]   _zz_io_p_95;
  reg        [47:0]   _zz_io_p_96;
  reg        [47:0]   _zz_io_p_97;
  reg        [47:0]   _zz_io_p_98;
  reg        [47:0]   _zz_io_p_99;
  reg        [47:0]   _zz_io_p_100;
  reg        [47:0]   _zz_io_p_101;
  reg        [47:0]   _zz_io_p_102;
  reg        [47:0]   _zz_io_p_103;
  reg        [47:0]   _zz_io_p_104;
  reg        [47:0]   _zz_io_p_105;
  reg        [47:0]   _zz_io_p_106;
  reg        [47:0]   _zz_io_p_107;
  reg        [47:0]   _zz_io_p_108;
  reg        [47:0]   _zz_io_p_109;
  reg        [47:0]   _zz_io_p_110;
  reg        [47:0]   _zz_io_p_111;
  reg        [47:0]   _zz_io_p_112;
  reg        [47:0]   _zz_io_p_113;
  reg        [47:0]   _zz_io_p_114;
  reg        [47:0]   _zz_io_p_115;
  reg        [47:0]   _zz_io_p_116;
  reg        [47:0]   _zz_io_p_117;
  reg        [47:0]   _zz_io_p_118;
  reg        [47:0]   _zz_io_p_119;
  reg        [47:0]   _zz_io_p_120;

  assign _zz_io_p_121 = _zz_io_p_75;
  assign _zz_io_p_122 = {_zz_io_p_65,{_zz_io_p_54,{_zz_io_p_42,{_zz_io_p_29,_zz_io_p_15}}}};
  KaratsubaCore_35 core (
    .io_a_0 (core_io_a_0[47:0]), //i
    .io_a_1 (core_io_a_1[47:0]), //i
    .io_a_2 (core_io_a_2[47:0]), //i
    .io_a_3 (core_io_a_3[47:0]), //i
    .io_a_4 (core_io_a_4[47:0]), //i
    .io_a_5 (core_io_a_5[47:0]), //i
    .io_a_6 (core_io_a_6[47:0]), //i
    .io_a_7 (core_io_a_7[47:0]), //i
    .io_b_0 (core_io_b_0[47:0]), //i
    .io_b_1 (core_io_b_1[47:0]), //i
    .io_b_2 (core_io_b_2[47:0]), //i
    .io_b_3 (core_io_b_3[47:0]), //i
    .io_b_4 (core_io_b_4[47:0]), //i
    .io_b_5 (core_io_b_5[47:0]), //i
    .io_b_6 (core_io_b_6[47:0]), //i
    .io_b_7 (core_io_b_7[47:0]), //i
    .io_p   (core_io_p[767:0] ), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  assign a = {7'd0, io_a};
  assign b = {7'd0, io_b};
  assign _zz_io_a_0 = a[335:0];
  assign core_io_a_0 = _zz_io_a_0[47 : 0];
  assign core_io_a_1 = _zz_io_a_0[95 : 48];
  assign core_io_a_2 = _zz_io_a_0[143 : 96];
  assign core_io_a_3 = _zz_io_a_0[191 : 144];
  assign core_io_a_4 = _zz_io_a_0[239 : 192];
  assign core_io_a_5 = _zz_io_a_0[287 : 240];
  assign core_io_a_6 = _zz_io_a_0[335 : 288];
  assign core_io_a_7 = (a >>> 336);
  assign _zz_io_b_0 = b[335:0];
  assign core_io_b_0 = _zz_io_b_0[47 : 0];
  assign core_io_b_1 = _zz_io_b_0[95 : 48];
  assign core_io_b_2 = _zz_io_b_0[143 : 96];
  assign core_io_b_3 = _zz_io_b_0[191 : 144];
  assign core_io_b_4 = _zz_io_b_0[239 : 192];
  assign core_io_b_5 = _zz_io_b_0[287 : 240];
  assign core_io_b_6 = _zz_io_b_0[335 : 288];
  assign core_io_b_7 = (b >>> 336);
  assign _zz_io_p = core_io_p[753:0];
  assign io_p = {_zz_io_p[753 : 720],{_zz_io_p_120,{_zz_io_p_119,{_zz_io_p_117,{_zz_io_p_114,{_zz_io_p_110,{_zz_io_p_105,{_zz_io_p_99,{_zz_io_p_92,{_zz_io_p_84,{_zz_io_p_121,_zz_io_p_122}}}}}}}}}}};
  always @(posedge clk) begin
    _zz_io_p_1 <= _zz_io_p[47 : 0];
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= _zz_io_p_2;
    _zz_io_p_4 <= _zz_io_p_3;
    _zz_io_p_5 <= _zz_io_p_4;
    _zz_io_p_6 <= _zz_io_p_5;
    _zz_io_p_7 <= _zz_io_p_6;
    _zz_io_p_8 <= _zz_io_p_7;
    _zz_io_p_9 <= _zz_io_p_8;
    _zz_io_p_10 <= _zz_io_p_9;
    _zz_io_p_11 <= _zz_io_p_10;
    _zz_io_p_12 <= _zz_io_p_11;
    _zz_io_p_13 <= _zz_io_p_12;
    _zz_io_p_14 <= _zz_io_p_13;
    _zz_io_p_15 <= _zz_io_p_14;
    _zz_io_p_16 <= _zz_io_p[95 : 48];
    _zz_io_p_17 <= _zz_io_p_16;
    _zz_io_p_18 <= _zz_io_p_17;
    _zz_io_p_19 <= _zz_io_p_18;
    _zz_io_p_20 <= _zz_io_p_19;
    _zz_io_p_21 <= _zz_io_p_20;
    _zz_io_p_22 <= _zz_io_p_21;
    _zz_io_p_23 <= _zz_io_p_22;
    _zz_io_p_24 <= _zz_io_p_23;
    _zz_io_p_25 <= _zz_io_p_24;
    _zz_io_p_26 <= _zz_io_p_25;
    _zz_io_p_27 <= _zz_io_p_26;
    _zz_io_p_28 <= _zz_io_p_27;
    _zz_io_p_29 <= _zz_io_p_28;
    _zz_io_p_30 <= _zz_io_p[143 : 96];
    _zz_io_p_31 <= _zz_io_p_30;
    _zz_io_p_32 <= _zz_io_p_31;
    _zz_io_p_33 <= _zz_io_p_32;
    _zz_io_p_34 <= _zz_io_p_33;
    _zz_io_p_35 <= _zz_io_p_34;
    _zz_io_p_36 <= _zz_io_p_35;
    _zz_io_p_37 <= _zz_io_p_36;
    _zz_io_p_38 <= _zz_io_p_37;
    _zz_io_p_39 <= _zz_io_p_38;
    _zz_io_p_40 <= _zz_io_p_39;
    _zz_io_p_41 <= _zz_io_p_40;
    _zz_io_p_42 <= _zz_io_p_41;
    _zz_io_p_43 <= _zz_io_p[191 : 144];
    _zz_io_p_44 <= _zz_io_p_43;
    _zz_io_p_45 <= _zz_io_p_44;
    _zz_io_p_46 <= _zz_io_p_45;
    _zz_io_p_47 <= _zz_io_p_46;
    _zz_io_p_48 <= _zz_io_p_47;
    _zz_io_p_49 <= _zz_io_p_48;
    _zz_io_p_50 <= _zz_io_p_49;
    _zz_io_p_51 <= _zz_io_p_50;
    _zz_io_p_52 <= _zz_io_p_51;
    _zz_io_p_53 <= _zz_io_p_52;
    _zz_io_p_54 <= _zz_io_p_53;
    _zz_io_p_55 <= _zz_io_p[239 : 192];
    _zz_io_p_56 <= _zz_io_p_55;
    _zz_io_p_57 <= _zz_io_p_56;
    _zz_io_p_58 <= _zz_io_p_57;
    _zz_io_p_59 <= _zz_io_p_58;
    _zz_io_p_60 <= _zz_io_p_59;
    _zz_io_p_61 <= _zz_io_p_60;
    _zz_io_p_62 <= _zz_io_p_61;
    _zz_io_p_63 <= _zz_io_p_62;
    _zz_io_p_64 <= _zz_io_p_63;
    _zz_io_p_65 <= _zz_io_p_64;
    _zz_io_p_66 <= _zz_io_p[287 : 240];
    _zz_io_p_67 <= _zz_io_p_66;
    _zz_io_p_68 <= _zz_io_p_67;
    _zz_io_p_69 <= _zz_io_p_68;
    _zz_io_p_70 <= _zz_io_p_69;
    _zz_io_p_71 <= _zz_io_p_70;
    _zz_io_p_72 <= _zz_io_p_71;
    _zz_io_p_73 <= _zz_io_p_72;
    _zz_io_p_74 <= _zz_io_p_73;
    _zz_io_p_75 <= _zz_io_p_74;
    _zz_io_p_76 <= _zz_io_p[335 : 288];
    _zz_io_p_77 <= _zz_io_p_76;
    _zz_io_p_78 <= _zz_io_p_77;
    _zz_io_p_79 <= _zz_io_p_78;
    _zz_io_p_80 <= _zz_io_p_79;
    _zz_io_p_81 <= _zz_io_p_80;
    _zz_io_p_82 <= _zz_io_p_81;
    _zz_io_p_83 <= _zz_io_p_82;
    _zz_io_p_84 <= _zz_io_p_83;
    _zz_io_p_85 <= _zz_io_p[383 : 336];
    _zz_io_p_86 <= _zz_io_p_85;
    _zz_io_p_87 <= _zz_io_p_86;
    _zz_io_p_88 <= _zz_io_p_87;
    _zz_io_p_89 <= _zz_io_p_88;
    _zz_io_p_90 <= _zz_io_p_89;
    _zz_io_p_91 <= _zz_io_p_90;
    _zz_io_p_92 <= _zz_io_p_91;
    _zz_io_p_93 <= _zz_io_p[431 : 384];
    _zz_io_p_94 <= _zz_io_p_93;
    _zz_io_p_95 <= _zz_io_p_94;
    _zz_io_p_96 <= _zz_io_p_95;
    _zz_io_p_97 <= _zz_io_p_96;
    _zz_io_p_98 <= _zz_io_p_97;
    _zz_io_p_99 <= _zz_io_p_98;
    _zz_io_p_100 <= _zz_io_p[479 : 432];
    _zz_io_p_101 <= _zz_io_p_100;
    _zz_io_p_102 <= _zz_io_p_101;
    _zz_io_p_103 <= _zz_io_p_102;
    _zz_io_p_104 <= _zz_io_p_103;
    _zz_io_p_105 <= _zz_io_p_104;
    _zz_io_p_106 <= _zz_io_p[527 : 480];
    _zz_io_p_107 <= _zz_io_p_106;
    _zz_io_p_108 <= _zz_io_p_107;
    _zz_io_p_109 <= _zz_io_p_108;
    _zz_io_p_110 <= _zz_io_p_109;
    _zz_io_p_111 <= _zz_io_p[575 : 528];
    _zz_io_p_112 <= _zz_io_p_111;
    _zz_io_p_113 <= _zz_io_p_112;
    _zz_io_p_114 <= _zz_io_p_113;
    _zz_io_p_115 <= _zz_io_p[623 : 576];
    _zz_io_p_116 <= _zz_io_p_115;
    _zz_io_p_117 <= _zz_io_p_116;
    _zz_io_p_118 <= _zz_io_p[671 : 624];
    _zz_io_p_119 <= _zz_io_p_118;
    _zz_io_p_120 <= _zz_io_p[719 : 672];
  end


endmodule

//ADD_11 replaced by ADD_5761

//ADD_10 replaced by ADD_5756

//ADD_9 replaced by ADD_5756

//ADD_8 replaced by ADD_5756

//ADD_7 replaced by ADD_5756

//ADD_6 replaced by ADD_5756

//BADD_37 replaced by BADD_1306

//ADD_17 replaced by ADD_167

//ADD_16 replaced by ADD_5756

//ADD_15 replaced by ADD_5756

//ADD_14 replaced by ADD_5756

//ADD_13 replaced by ADD_5756

//ADD_12 replaced by ADD_5756

//BADD_38 replaced by BADD_1306

//ADD_23 replaced by ADD_167

//ADD_22 replaced by ADD_5756

//ADD_21 replaced by ADD_5756

//ADD_20 replaced by ADD_5756

//ADD_19 replaced by ADD_5756

//ADD_18 replaced by ADD_5756

//BADD_39 replaced by BADD_1306

//ADD_29 replaced by ADD_167

//ADD_28 replaced by ADD_5756

//ADD_27 replaced by ADD_5756

//ADD_26 replaced by ADD_5756

//ADD_25 replaced by ADD_5756

//ADD_24 replaced by ADD_5756

//BADD_40 replaced by BADD_1306

//ADD_35 replaced by ADD_167

//ADD_34 replaced by ADD_5756

//ADD_33 replaced by ADD_5756

//ADD_32 replaced by ADD_5756

//ADD_31 replaced by ADD_5756

//ADD_30 replaced by ADD_5756

//BADD_41 replaced by BADD_619

//ADD_41 replaced by ADD_167

//ADD_40 replaced by ADD_5756

//ADD_39 replaced by ADD_5756

//ADD_38 replaced by ADD_5756

//ADD_37 replaced by ADD_5756

//ADD_36 replaced by ADD_5756

//BADD_42 replaced by BADD_619

//ADD_47 replaced by ADD_167

//ADD_46 replaced by ADD_5756

//ADD_45 replaced by ADD_5756

//ADD_44 replaced by ADD_5756

//ADD_43 replaced by ADD_5756

//ADD_42 replaced by ADD_5756

//BADD_43 replaced by BADD_619

//ADD_53 replaced by ADD_167

//ADD_52 replaced by ADD_5756

//ADD_51 replaced by ADD_5756

//ADD_50 replaced by ADD_5756

//ADD_49 replaced by ADD_5756

//ADD_48 replaced by ADD_5756

//BADD_44 replaced by BADD_619

//ADD_59 replaced by ADD_167

//ADD_58 replaced by ADD_5756

//ADD_57 replaced by ADD_5756

//ADD_56 replaced by ADD_5756

//ADD_55 replaced by ADD_5756

//ADD_54 replaced by ADD_5756

//FineReduction_36 replaced by FineReduction_53

//BADD_45 replaced by BADD_1124

//ADD_65 replaced by ADD_4223

//ADD_64 replaced by ADD_5756

//ADD_63 replaced by ADD_5756

//ADD_62 replaced by ADD_5756

//ADD_61 replaced by ADD_5756

//ADD_60 replaced by ADD_5756

//BADD_107 replaced by BADD_1186

//BADD_106 replaced by BADD_1185

//BADD_105 replaced by BADD_1184

//BADD_104 replaced by BADD_1183

//BADD_103 replaced by BADD_1182

//BADD_102 replaced by BADD_1181

//BADD_101 replaced by BADD_1180

//BADD_100 replaced by BADD_1179

//BADD_99 replaced by BADD_1178

//BADD_98 replaced by BADD_1177

//BADD_97 replaced by BADD_1176

//BADD_96 replaced by BADD_1175

//BADD_95 replaced by BADD_1174

//BADD_94 replaced by BADD_1173

//BADD_93 replaced by BADD_1172

//BADD_92 replaced by BADD_1171

//BADD_91 replaced by BADD_1170

//BADD_90 replaced by BADD_1169

//BADD_89 replaced by BADD_1168

//BADD_88 replaced by BADD_1167

//BADD_87 replaced by BADD_1166

//BADD_86 replaced by BADD_1165

//BADD_85 replaced by BADD_1164

//BADD_84 replaced by BADD_1163

//BADD_83 replaced by BADD_1162

//BADD_82 replaced by BADD_1161

//BADD_81 replaced by BADD_1160

//BADD_80 replaced by BADD_1159

//BADD_79 replaced by BADD_1158

//BADD_78 replaced by BADD_1157

//BADD_77 replaced by BADD_1156

//BADD_76 replaced by BADD_1155

//BADD_75 replaced by BADD_1154

//BADD_74 replaced by BADD_1153

//BADD_73 replaced by BADD_1152

//BADD_72 replaced by BADD_1151

//BADD_71 replaced by BADD_1150

//BADD_70 replaced by BADD_1149

//BADD_69 replaced by BADD_1148

//BADD_68 replaced by BADD_1147

//BADD_67 replaced by BADD_1146

//BADD_66 replaced by BADD_1145

//BADD_65 replaced by BADD_1144

//BADD_64 replaced by BADD_1143

//BADD_63 replaced by BADD_1142

//BADD_62 replaced by BADD_1141

//BADD_61 replaced by BADD_1140

//BADD_60 replaced by BADD_1139

//BADD_59 replaced by BADD_1138

//BADD_58 replaced by BADD_1137

//BADD_57 replaced by BADD_1136

//BADD_56 replaced by BADD_1135

//BADD_55 replaced by BADD_1134

//BADD_54 replaced by BADD_1133

//BADD_53 replaced by BADD_1132

//BADD_52 replaced by BADD_1131

//BADD_51 replaced by BADD_1130

//BADD_50 replaced by BADD_1129

//BADD_49 replaced by BADD_1128

//BADD_48 replaced by BADD_1127

//BADD_47 replaced by BADD_1126

//BADD_46 replaced by BADD_1125

//KaratsubaCore replaced by KaratsubaCore_35

//KaratsubaCore_1 replaced by KaratsubaCore_35

//FineReduction_37 replaced by FineReduction_53

//BADD_108 replaced by BADD_1124

//ADD_71 replaced by ADD_4223

//ADD_70 replaced by ADD_5756

//ADD_69 replaced by ADD_5756

//ADD_68 replaced by ADD_5756

//ADD_67 replaced by ADD_5756

//ADD_66 replaced by ADD_5756

//BADD_170 replaced by BADD_1186

//BADD_169 replaced by BADD_1185

//BADD_168 replaced by BADD_1184

//BADD_167 replaced by BADD_1183

//BADD_166 replaced by BADD_1182

//BADD_165 replaced by BADD_1181

//BADD_164 replaced by BADD_1180

//BADD_163 replaced by BADD_1179

//BADD_162 replaced by BADD_1178

//BADD_161 replaced by BADD_1177

//BADD_160 replaced by BADD_1176

//BADD_159 replaced by BADD_1175

//BADD_158 replaced by BADD_1174

//BADD_157 replaced by BADD_1173

//BADD_156 replaced by BADD_1172

//BADD_155 replaced by BADD_1171

//BADD_154 replaced by BADD_1170

//BADD_153 replaced by BADD_1169

//BADD_152 replaced by BADD_1168

//BADD_151 replaced by BADD_1167

//BADD_150 replaced by BADD_1166

//BADD_149 replaced by BADD_1165

//BADD_148 replaced by BADD_1164

//BADD_147 replaced by BADD_1163

//BADD_146 replaced by BADD_1162

//BADD_145 replaced by BADD_1161

//BADD_144 replaced by BADD_1160

//BADD_143 replaced by BADD_1159

//BADD_142 replaced by BADD_1158

//BADD_141 replaced by BADD_1157

//BADD_140 replaced by BADD_1156

//BADD_139 replaced by BADD_1155

//BADD_138 replaced by BADD_1154

//BADD_137 replaced by BADD_1153

//BADD_136 replaced by BADD_1152

//BADD_135 replaced by BADD_1151

//BADD_134 replaced by BADD_1150

//BADD_133 replaced by BADD_1149

//BADD_132 replaced by BADD_1148

//BADD_131 replaced by BADD_1147

//BADD_130 replaced by BADD_1146

//BADD_129 replaced by BADD_1145

//BADD_128 replaced by BADD_1144

//BADD_127 replaced by BADD_1143

//BADD_126 replaced by BADD_1142

//BADD_125 replaced by BADD_1141

//BADD_124 replaced by BADD_1140

//BADD_123 replaced by BADD_1139

//BADD_122 replaced by BADD_1138

//BADD_121 replaced by BADD_1137

//BADD_120 replaced by BADD_1136

//BADD_119 replaced by BADD_1135

//BADD_118 replaced by BADD_1134

//BADD_117 replaced by BADD_1133

//BADD_116 replaced by BADD_1132

//BADD_115 replaced by BADD_1131

//BADD_114 replaced by BADD_1130

//BADD_113 replaced by BADD_1129

//BADD_112 replaced by BADD_1128

//BADD_111 replaced by BADD_1127

//BADD_110 replaced by BADD_1126

//BADD_109 replaced by BADD_1125

//KaratsubaCore_2 replaced by KaratsubaCore_35

//KaratsubaCore_3 replaced by KaratsubaCore_35

//FineReduction_38 replaced by FineReduction_53

//BADD_171 replaced by BADD_1124

//ADD_77 replaced by ADD_4223

//ADD_76 replaced by ADD_5756

//ADD_75 replaced by ADD_5756

//ADD_74 replaced by ADD_5756

//ADD_73 replaced by ADD_5756

//ADD_72 replaced by ADD_5756

//BADD_233 replaced by BADD_1186

//BADD_232 replaced by BADD_1185

//BADD_231 replaced by BADD_1184

//BADD_230 replaced by BADD_1183

//BADD_229 replaced by BADD_1182

//BADD_228 replaced by BADD_1181

//BADD_227 replaced by BADD_1180

//BADD_226 replaced by BADD_1179

//BADD_225 replaced by BADD_1178

//BADD_224 replaced by BADD_1177

//BADD_223 replaced by BADD_1176

//BADD_222 replaced by BADD_1175

//BADD_221 replaced by BADD_1174

//BADD_220 replaced by BADD_1173

//BADD_219 replaced by BADD_1172

//BADD_218 replaced by BADD_1171

//BADD_217 replaced by BADD_1170

//BADD_216 replaced by BADD_1169

//BADD_215 replaced by BADD_1168

//BADD_214 replaced by BADD_1167

//BADD_213 replaced by BADD_1166

//BADD_212 replaced by BADD_1165

//BADD_211 replaced by BADD_1164

//BADD_210 replaced by BADD_1163

//BADD_209 replaced by BADD_1162

//BADD_208 replaced by BADD_1161

//BADD_207 replaced by BADD_1160

//BADD_206 replaced by BADD_1159

//BADD_205 replaced by BADD_1158

//BADD_204 replaced by BADD_1157

//BADD_203 replaced by BADD_1156

//BADD_202 replaced by BADD_1155

//BADD_201 replaced by BADD_1154

//BADD_200 replaced by BADD_1153

//BADD_199 replaced by BADD_1152

//BADD_198 replaced by BADD_1151

//BADD_197 replaced by BADD_1150

//BADD_196 replaced by BADD_1149

//BADD_195 replaced by BADD_1148

//BADD_194 replaced by BADD_1147

//BADD_193 replaced by BADD_1146

//BADD_192 replaced by BADD_1145

//BADD_191 replaced by BADD_1144

//BADD_190 replaced by BADD_1143

//BADD_189 replaced by BADD_1142

//BADD_188 replaced by BADD_1141

//BADD_187 replaced by BADD_1140

//BADD_186 replaced by BADD_1139

//BADD_185 replaced by BADD_1138

//BADD_184 replaced by BADD_1137

//BADD_183 replaced by BADD_1136

//BADD_182 replaced by BADD_1135

//BADD_181 replaced by BADD_1134

//BADD_180 replaced by BADD_1133

//BADD_179 replaced by BADD_1132

//BADD_178 replaced by BADD_1131

//BADD_177 replaced by BADD_1130

//BADD_176 replaced by BADD_1129

//BADD_175 replaced by BADD_1128

//BADD_174 replaced by BADD_1127

//BADD_173 replaced by BADD_1126

//BADD_172 replaced by BADD_1125

//KaratsubaCore_4 replaced by KaratsubaCore_35

//KaratsubaCore_5 replaced by KaratsubaCore_35

//FineReduction_39 replaced by FineReduction_53

//BADD_234 replaced by BADD_1124

//ADD_83 replaced by ADD_4223

//ADD_82 replaced by ADD_5756

//ADD_81 replaced by ADD_5756

//ADD_80 replaced by ADD_5756

//ADD_79 replaced by ADD_5756

//ADD_78 replaced by ADD_5756

//BADD_296 replaced by BADD_1186

//BADD_295 replaced by BADD_1185

//BADD_294 replaced by BADD_1184

//BADD_293 replaced by BADD_1183

//BADD_292 replaced by BADD_1182

//BADD_291 replaced by BADD_1181

//BADD_290 replaced by BADD_1180

//BADD_289 replaced by BADD_1179

//BADD_288 replaced by BADD_1178

//BADD_287 replaced by BADD_1177

//BADD_286 replaced by BADD_1176

//BADD_285 replaced by BADD_1175

//BADD_284 replaced by BADD_1174

//BADD_283 replaced by BADD_1173

//BADD_282 replaced by BADD_1172

//BADD_281 replaced by BADD_1171

//BADD_280 replaced by BADD_1170

//BADD_279 replaced by BADD_1169

//BADD_278 replaced by BADD_1168

//BADD_277 replaced by BADD_1167

//BADD_276 replaced by BADD_1166

//BADD_275 replaced by BADD_1165

//BADD_274 replaced by BADD_1164

//BADD_273 replaced by BADD_1163

//BADD_272 replaced by BADD_1162

//BADD_271 replaced by BADD_1161

//BADD_270 replaced by BADD_1160

//BADD_269 replaced by BADD_1159

//BADD_268 replaced by BADD_1158

//BADD_267 replaced by BADD_1157

//BADD_266 replaced by BADD_1156

//BADD_265 replaced by BADD_1155

//BADD_264 replaced by BADD_1154

//BADD_263 replaced by BADD_1153

//BADD_262 replaced by BADD_1152

//BADD_261 replaced by BADD_1151

//BADD_260 replaced by BADD_1150

//BADD_259 replaced by BADD_1149

//BADD_258 replaced by BADD_1148

//BADD_257 replaced by BADD_1147

//BADD_256 replaced by BADD_1146

//BADD_255 replaced by BADD_1145

//BADD_254 replaced by BADD_1144

//BADD_253 replaced by BADD_1143

//BADD_252 replaced by BADD_1142

//BADD_251 replaced by BADD_1141

//BADD_250 replaced by BADD_1140

//BADD_249 replaced by BADD_1139

//BADD_248 replaced by BADD_1138

//BADD_247 replaced by BADD_1137

//BADD_246 replaced by BADD_1136

//BADD_245 replaced by BADD_1135

//BADD_244 replaced by BADD_1134

//BADD_243 replaced by BADD_1133

//BADD_242 replaced by BADD_1132

//BADD_241 replaced by BADD_1131

//BADD_240 replaced by BADD_1130

//BADD_239 replaced by BADD_1129

//BADD_238 replaced by BADD_1128

//BADD_237 replaced by BADD_1127

//BADD_236 replaced by BADD_1126

//BADD_235 replaced by BADD_1125

//KaratsubaCore_6 replaced by KaratsubaCore_35

//KaratsubaCore_7 replaced by KaratsubaCore_35

//FineReduction_40 replaced by FineReduction_53

//BADD_297 replaced by BADD_1124

//ADD_89 replaced by ADD_4223

//ADD_88 replaced by ADD_5756

//ADD_87 replaced by ADD_5756

//ADD_86 replaced by ADD_5756

//ADD_85 replaced by ADD_5756

//ADD_84 replaced by ADD_5756

//BADD_359 replaced by BADD_1186

//BADD_358 replaced by BADD_1185

//BADD_357 replaced by BADD_1184

//BADD_356 replaced by BADD_1183

//BADD_355 replaced by BADD_1182

//BADD_354 replaced by BADD_1181

//BADD_353 replaced by BADD_1180

//BADD_352 replaced by BADD_1179

//BADD_351 replaced by BADD_1178

//BADD_350 replaced by BADD_1177

//BADD_349 replaced by BADD_1176

//BADD_348 replaced by BADD_1175

//BADD_347 replaced by BADD_1174

//BADD_346 replaced by BADD_1173

//BADD_345 replaced by BADD_1172

//BADD_344 replaced by BADD_1171

//BADD_343 replaced by BADD_1170

//BADD_342 replaced by BADD_1169

//BADD_341 replaced by BADD_1168

//BADD_340 replaced by BADD_1167

//BADD_339 replaced by BADD_1166

//BADD_338 replaced by BADD_1165

//BADD_337 replaced by BADD_1164

//BADD_336 replaced by BADD_1163

//BADD_335 replaced by BADD_1162

//BADD_334 replaced by BADD_1161

//BADD_333 replaced by BADD_1160

//BADD_332 replaced by BADD_1159

//BADD_331 replaced by BADD_1158

//BADD_330 replaced by BADD_1157

//BADD_329 replaced by BADD_1156

//BADD_328 replaced by BADD_1155

//BADD_327 replaced by BADD_1154

//BADD_326 replaced by BADD_1153

//BADD_325 replaced by BADD_1152

//BADD_324 replaced by BADD_1151

//BADD_323 replaced by BADD_1150

//BADD_322 replaced by BADD_1149

//BADD_321 replaced by BADD_1148

//BADD_320 replaced by BADD_1147

//BADD_319 replaced by BADD_1146

//BADD_318 replaced by BADD_1145

//BADD_317 replaced by BADD_1144

//BADD_316 replaced by BADD_1143

//BADD_315 replaced by BADD_1142

//BADD_314 replaced by BADD_1141

//BADD_313 replaced by BADD_1140

//BADD_312 replaced by BADD_1139

//BADD_311 replaced by BADD_1138

//BADD_310 replaced by BADD_1137

//BADD_309 replaced by BADD_1136

//BADD_308 replaced by BADD_1135

//BADD_307 replaced by BADD_1134

//BADD_306 replaced by BADD_1133

//BADD_305 replaced by BADD_1132

//BADD_304 replaced by BADD_1131

//BADD_303 replaced by BADD_1130

//BADD_302 replaced by BADD_1129

//BADD_301 replaced by BADD_1128

//BADD_300 replaced by BADD_1127

//BADD_299 replaced by BADD_1126

//BADD_298 replaced by BADD_1125

//KaratsubaCore_8 replaced by KaratsubaCore_35

//KaratsubaCore_9 replaced by KaratsubaCore_35

//FineReduction_41 replaced by FineReduction_53

//BADD_360 replaced by BADD_1124

//ADD_95 replaced by ADD_4223

//ADD_94 replaced by ADD_5756

//ADD_93 replaced by ADD_5756

//ADD_92 replaced by ADD_5756

//ADD_91 replaced by ADD_5756

//ADD_90 replaced by ADD_5756

//BADD_422 replaced by BADD_1186

//BADD_421 replaced by BADD_1185

//BADD_420 replaced by BADD_1184

//BADD_419 replaced by BADD_1183

//BADD_418 replaced by BADD_1182

//BADD_417 replaced by BADD_1181

//BADD_416 replaced by BADD_1180

//BADD_415 replaced by BADD_1179

//BADD_414 replaced by BADD_1178

//BADD_413 replaced by BADD_1177

//BADD_412 replaced by BADD_1176

//BADD_411 replaced by BADD_1175

//BADD_410 replaced by BADD_1174

//BADD_409 replaced by BADD_1173

//BADD_408 replaced by BADD_1172

//BADD_407 replaced by BADD_1171

//BADD_406 replaced by BADD_1170

//BADD_405 replaced by BADD_1169

//BADD_404 replaced by BADD_1168

//BADD_403 replaced by BADD_1167

//BADD_402 replaced by BADD_1166

//BADD_401 replaced by BADD_1165

//BADD_400 replaced by BADD_1164

//BADD_399 replaced by BADD_1163

//BADD_398 replaced by BADD_1162

//BADD_397 replaced by BADD_1161

//BADD_396 replaced by BADD_1160

//BADD_395 replaced by BADD_1159

//BADD_394 replaced by BADD_1158

//BADD_393 replaced by BADD_1157

//BADD_392 replaced by BADD_1156

//BADD_391 replaced by BADD_1155

//BADD_390 replaced by BADD_1154

//BADD_389 replaced by BADD_1153

//BADD_388 replaced by BADD_1152

//BADD_387 replaced by BADD_1151

//BADD_386 replaced by BADD_1150

//BADD_385 replaced by BADD_1149

//BADD_384 replaced by BADD_1148

//BADD_383 replaced by BADD_1147

//BADD_382 replaced by BADD_1146

//BADD_381 replaced by BADD_1145

//BADD_380 replaced by BADD_1144

//BADD_379 replaced by BADD_1143

//BADD_378 replaced by BADD_1142

//BADD_377 replaced by BADD_1141

//BADD_376 replaced by BADD_1140

//BADD_375 replaced by BADD_1139

//BADD_374 replaced by BADD_1138

//BADD_373 replaced by BADD_1137

//BADD_372 replaced by BADD_1136

//BADD_371 replaced by BADD_1135

//BADD_370 replaced by BADD_1134

//BADD_369 replaced by BADD_1133

//BADD_368 replaced by BADD_1132

//BADD_367 replaced by BADD_1131

//BADD_366 replaced by BADD_1130

//BADD_365 replaced by BADD_1129

//BADD_364 replaced by BADD_1128

//BADD_363 replaced by BADD_1127

//BADD_362 replaced by BADD_1126

//BADD_361 replaced by BADD_1125

//KaratsubaCore_10 replaced by KaratsubaCore_35

//KaratsubaCore_11 replaced by KaratsubaCore_35

//FineReduction_42 replaced by FineReduction_53

//BADD_423 replaced by BADD_1124

//ADD_101 replaced by ADD_4223

//ADD_100 replaced by ADD_5756

//ADD_99 replaced by ADD_5756

//ADD_98 replaced by ADD_5756

//ADD_97 replaced by ADD_5756

//ADD_96 replaced by ADD_5756

//BADD_485 replaced by BADD_1186

//BADD_484 replaced by BADD_1185

//BADD_483 replaced by BADD_1184

//BADD_482 replaced by BADD_1183

//BADD_481 replaced by BADD_1182

//BADD_480 replaced by BADD_1181

//BADD_479 replaced by BADD_1180

//BADD_478 replaced by BADD_1179

//BADD_477 replaced by BADD_1178

//BADD_476 replaced by BADD_1177

//BADD_475 replaced by BADD_1176

//BADD_474 replaced by BADD_1175

//BADD_473 replaced by BADD_1174

//BADD_472 replaced by BADD_1173

//BADD_471 replaced by BADD_1172

//BADD_470 replaced by BADD_1171

//BADD_469 replaced by BADD_1170

//BADD_468 replaced by BADD_1169

//BADD_467 replaced by BADD_1168

//BADD_466 replaced by BADD_1167

//BADD_465 replaced by BADD_1166

//BADD_464 replaced by BADD_1165

//BADD_463 replaced by BADD_1164

//BADD_462 replaced by BADD_1163

//BADD_461 replaced by BADD_1162

//BADD_460 replaced by BADD_1161

//BADD_459 replaced by BADD_1160

//BADD_458 replaced by BADD_1159

//BADD_457 replaced by BADD_1158

//BADD_456 replaced by BADD_1157

//BADD_455 replaced by BADD_1156

//BADD_454 replaced by BADD_1155

//BADD_453 replaced by BADD_1154

//BADD_452 replaced by BADD_1153

//BADD_451 replaced by BADD_1152

//BADD_450 replaced by BADD_1151

//BADD_449 replaced by BADD_1150

//BADD_448 replaced by BADD_1149

//BADD_447 replaced by BADD_1148

//BADD_446 replaced by BADD_1147

//BADD_445 replaced by BADD_1146

//BADD_444 replaced by BADD_1145

//BADD_443 replaced by BADD_1144

//BADD_442 replaced by BADD_1143

//BADD_441 replaced by BADD_1142

//BADD_440 replaced by BADD_1141

//BADD_439 replaced by BADD_1140

//BADD_438 replaced by BADD_1139

//BADD_437 replaced by BADD_1138

//BADD_436 replaced by BADD_1137

//BADD_435 replaced by BADD_1136

//BADD_434 replaced by BADD_1135

//BADD_433 replaced by BADD_1134

//BADD_432 replaced by BADD_1133

//BADD_431 replaced by BADD_1132

//BADD_430 replaced by BADD_1131

//BADD_429 replaced by BADD_1130

//BADD_428 replaced by BADD_1129

//BADD_427 replaced by BADD_1128

//BADD_426 replaced by BADD_1127

//BADD_425 replaced by BADD_1126

//BADD_424 replaced by BADD_1125

//KaratsubaCore_12 replaced by KaratsubaCore_35

//KaratsubaCore_13 replaced by KaratsubaCore_35

//FineReduction_43 replaced by FineReduction_53

//BADD_486 replaced by BADD_1124

//ADD_107 replaced by ADD_4223

//ADD_106 replaced by ADD_5756

//ADD_105 replaced by ADD_5756

//ADD_104 replaced by ADD_5756

//ADD_103 replaced by ADD_5756

//ADD_102 replaced by ADD_5756

//BADD_548 replaced by BADD_1186

//BADD_547 replaced by BADD_1185

//BADD_546 replaced by BADD_1184

//BADD_545 replaced by BADD_1183

//BADD_544 replaced by BADD_1182

//BADD_543 replaced by BADD_1181

//BADD_542 replaced by BADD_1180

//BADD_541 replaced by BADD_1179

//BADD_540 replaced by BADD_1178

//BADD_539 replaced by BADD_1177

//BADD_538 replaced by BADD_1176

//BADD_537 replaced by BADD_1175

//BADD_536 replaced by BADD_1174

//BADD_535 replaced by BADD_1173

//BADD_534 replaced by BADD_1172

//BADD_533 replaced by BADD_1171

//BADD_532 replaced by BADD_1170

//BADD_531 replaced by BADD_1169

//BADD_530 replaced by BADD_1168

//BADD_529 replaced by BADD_1167

//BADD_528 replaced by BADD_1166

//BADD_527 replaced by BADD_1165

//BADD_526 replaced by BADD_1164

//BADD_525 replaced by BADD_1163

//BADD_524 replaced by BADD_1162

//BADD_523 replaced by BADD_1161

//BADD_522 replaced by BADD_1160

//BADD_521 replaced by BADD_1159

//BADD_520 replaced by BADD_1158

//BADD_519 replaced by BADD_1157

//BADD_518 replaced by BADD_1156

//BADD_517 replaced by BADD_1155

//BADD_516 replaced by BADD_1154

//BADD_515 replaced by BADD_1153

//BADD_514 replaced by BADD_1152

//BADD_513 replaced by BADD_1151

//BADD_512 replaced by BADD_1150

//BADD_511 replaced by BADD_1149

//BADD_510 replaced by BADD_1148

//BADD_509 replaced by BADD_1147

//BADD_508 replaced by BADD_1146

//BADD_507 replaced by BADD_1145

//BADD_506 replaced by BADD_1144

//BADD_505 replaced by BADD_1143

//BADD_504 replaced by BADD_1142

//BADD_503 replaced by BADD_1141

//BADD_502 replaced by BADD_1140

//BADD_501 replaced by BADD_1139

//BADD_500 replaced by BADD_1138

//BADD_499 replaced by BADD_1137

//BADD_498 replaced by BADD_1136

//BADD_497 replaced by BADD_1135

//BADD_496 replaced by BADD_1134

//BADD_495 replaced by BADD_1133

//BADD_494 replaced by BADD_1132

//BADD_493 replaced by BADD_1131

//BADD_492 replaced by BADD_1130

//BADD_491 replaced by BADD_1129

//BADD_490 replaced by BADD_1128

//BADD_489 replaced by BADD_1127

//BADD_488 replaced by BADD_1126

//BADD_487 replaced by BADD_1125

//KaratsubaCore_14 replaced by KaratsubaCore_35

//KaratsubaCore_15 replaced by KaratsubaCore_35

//FineReduction_44 replaced by FineReduction_53

//BADD_549 replaced by BADD_1124

//ADD_113 replaced by ADD_4223

//ADD_112 replaced by ADD_5756

//ADD_111 replaced by ADD_5756

//ADD_110 replaced by ADD_5756

//ADD_109 replaced by ADD_5756

//ADD_108 replaced by ADD_5756

//BADD_611 replaced by BADD_1186

//BADD_610 replaced by BADD_1185

//BADD_609 replaced by BADD_1184

//BADD_608 replaced by BADD_1183

//BADD_607 replaced by BADD_1182

//BADD_606 replaced by BADD_1181

//BADD_605 replaced by BADD_1180

//BADD_604 replaced by BADD_1179

//BADD_603 replaced by BADD_1178

//BADD_602 replaced by BADD_1177

//BADD_601 replaced by BADD_1176

//BADD_600 replaced by BADD_1175

//BADD_599 replaced by BADD_1174

//BADD_598 replaced by BADD_1173

//BADD_597 replaced by BADD_1172

//BADD_596 replaced by BADD_1171

//BADD_595 replaced by BADD_1170

//BADD_594 replaced by BADD_1169

//BADD_593 replaced by BADD_1168

//BADD_592 replaced by BADD_1167

//BADD_591 replaced by BADD_1166

//BADD_590 replaced by BADD_1165

//BADD_589 replaced by BADD_1164

//BADD_588 replaced by BADD_1163

//BADD_587 replaced by BADD_1162

//BADD_586 replaced by BADD_1161

//BADD_585 replaced by BADD_1160

//BADD_584 replaced by BADD_1159

//BADD_583 replaced by BADD_1158

//BADD_582 replaced by BADD_1157

//BADD_581 replaced by BADD_1156

//BADD_580 replaced by BADD_1155

//BADD_579 replaced by BADD_1154

//BADD_578 replaced by BADD_1153

//BADD_577 replaced by BADD_1152

//BADD_576 replaced by BADD_1151

//BADD_575 replaced by BADD_1150

//BADD_574 replaced by BADD_1149

//BADD_573 replaced by BADD_1148

//BADD_572 replaced by BADD_1147

//BADD_571 replaced by BADD_1146

//BADD_570 replaced by BADD_1145

//BADD_569 replaced by BADD_1144

//BADD_568 replaced by BADD_1143

//BADD_567 replaced by BADD_1142

//BADD_566 replaced by BADD_1141

//BADD_565 replaced by BADD_1140

//BADD_564 replaced by BADD_1139

//BADD_563 replaced by BADD_1138

//BADD_562 replaced by BADD_1137

//BADD_561 replaced by BADD_1136

//BADD_560 replaced by BADD_1135

//BADD_559 replaced by BADD_1134

//BADD_558 replaced by BADD_1133

//BADD_557 replaced by BADD_1132

//BADD_556 replaced by BADD_1131

//BADD_555 replaced by BADD_1130

//BADD_554 replaced by BADD_1129

//BADD_553 replaced by BADD_1128

//BADD_552 replaced by BADD_1127

//BADD_551 replaced by BADD_1126

//BADD_550 replaced by BADD_1125

//KaratsubaCore_16 replaced by KaratsubaCore_35

//KaratsubaCore_17 replaced by KaratsubaCore_35

//ADD_119 replaced by ADD_5761

//ADD_118 replaced by ADD_5756

//ADD_117 replaced by ADD_5756

//ADD_116 replaced by ADD_5756

//ADD_115 replaced by ADD_5756

//ADD_114 replaced by ADD_5756

//BADD_612 replaced by BADD_1306

//ADD_125 replaced by ADD_167

//ADD_124 replaced by ADD_5756

//ADD_123 replaced by ADD_5756

//ADD_122 replaced by ADD_5756

//ADD_121 replaced by ADD_5756

//ADD_120 replaced by ADD_5756

//BADD_613 replaced by BADD_1306

//ADD_131 replaced by ADD_167

//ADD_130 replaced by ADD_5756

//ADD_129 replaced by ADD_5756

//ADD_128 replaced by ADD_5756

//ADD_127 replaced by ADD_5756

//ADD_126 replaced by ADD_5756

//BADD_614 replaced by BADD_1306

//ADD_137 replaced by ADD_167

//ADD_136 replaced by ADD_5756

//ADD_135 replaced by ADD_5756

//ADD_134 replaced by ADD_5756

//ADD_133 replaced by ADD_5756

//ADD_132 replaced by ADD_5756

//BADD_615 replaced by BADD_1306

//ADD_143 replaced by ADD_167

//ADD_142 replaced by ADD_5756

//ADD_141 replaced by ADD_5756

//ADD_140 replaced by ADD_5756

//ADD_139 replaced by ADD_5756

//ADD_138 replaced by ADD_5756

//BADD_616 replaced by BADD_619

//ADD_149 replaced by ADD_167

//ADD_148 replaced by ADD_5756

//ADD_147 replaced by ADD_5756

//ADD_146 replaced by ADD_5756

//ADD_145 replaced by ADD_5756

//ADD_144 replaced by ADD_5756

//BADD_617 replaced by BADD_619

//ADD_155 replaced by ADD_167

//ADD_154 replaced by ADD_5756

//ADD_153 replaced by ADD_5756

//ADD_152 replaced by ADD_5756

//ADD_151 replaced by ADD_5756

//ADD_150 replaced by ADD_5756

//BADD_618 replaced by BADD_619

//ADD_161 replaced by ADD_167

//ADD_160 replaced by ADD_5756

//ADD_159 replaced by ADD_5756

//ADD_158 replaced by ADD_5756

//ADD_157 replaced by ADD_5756

//ADD_156 replaced by ADD_5756

module BADD_619 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  input               io_c,
  output     [378:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [57:0]   adder_adds_5_io_A_0;
  wire       [57:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [58:0]   adder_adds_5_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  reg        [57:0]   _zz_io_s_21;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_5761 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[57:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[57:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[58:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = io_a[127 : 64];
  assign adder_adds_2_io_A_0 = io_a[191 : 128];
  assign adder_adds_3_io_A_0 = io_a[255 : 192];
  assign adder_adds_4_io_A_0 = io_a[319 : 256];
  assign adder_adds_5_io_A_0 = io_a[377 : 320];
  assign adder_adds_0_io_A_1 = (~ io_b[63 : 0]);
  assign adder_adds_1_io_A_1 = (~ io_b[127 : 64]);
  assign adder_adds_2_io_A_1 = (~ io_b[191 : 128]);
  assign adder_adds_3_io_A_1 = (~ io_b[255 : 192]);
  assign adder_adds_4_io_A_1 = (~ io_b[319 : 256]);
  assign adder_adds_5_io_A_1 = (~ io_b[377 : 320]);
  assign io_s = {_zz_io_s,{_zz_io_s_21,{_zz_io_s_20,{_zz_io_s_18,{_zz_io_s_15,{_zz_io_s_11,_zz_io_s_6}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= (! adder_adds_5_io_S[58]);
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_8 <= _zz_io_s_7;
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_21 <= adder_adds_5_io_S[57 : 0];
  end


endmodule

module ADD_167 (
  input      [56:0]   io_A_0,
  input      [56:0]   io_A_1,
  input               io_CIN,
  output     [57:0]   io_S
);

  wire       [57:0]   _zz_io_S;
  wire       [57:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {57'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_166 replaced by ADD_5756

//ADD_165 replaced by ADD_5756

//ADD_164 replaced by ADD_5756

//ADD_163 replaced by ADD_5756

//ADD_162 replaced by ADD_5756

//FineReduction_45 replaced by FineReduction_53

//BADD_620 replaced by BADD_1124

//ADD_173 replaced by ADD_4223

//ADD_172 replaced by ADD_5756

//ADD_171 replaced by ADD_5756

//ADD_170 replaced by ADD_5756

//ADD_169 replaced by ADD_5756

//ADD_168 replaced by ADD_5756

//BADD_682 replaced by BADD_1186

//BADD_681 replaced by BADD_1185

//BADD_680 replaced by BADD_1184

//BADD_679 replaced by BADD_1183

//BADD_678 replaced by BADD_1182

//BADD_677 replaced by BADD_1181

//BADD_676 replaced by BADD_1180

//BADD_675 replaced by BADD_1179

//BADD_674 replaced by BADD_1178

//BADD_673 replaced by BADD_1177

//BADD_672 replaced by BADD_1176

//BADD_671 replaced by BADD_1175

//BADD_670 replaced by BADD_1174

//BADD_669 replaced by BADD_1173

//BADD_668 replaced by BADD_1172

//BADD_667 replaced by BADD_1171

//BADD_666 replaced by BADD_1170

//BADD_665 replaced by BADD_1169

//BADD_664 replaced by BADD_1168

//BADD_663 replaced by BADD_1167

//BADD_662 replaced by BADD_1166

//BADD_661 replaced by BADD_1165

//BADD_660 replaced by BADD_1164

//BADD_659 replaced by BADD_1163

//BADD_658 replaced by BADD_1162

//BADD_657 replaced by BADD_1161

//BADD_656 replaced by BADD_1160

//BADD_655 replaced by BADD_1159

//BADD_654 replaced by BADD_1158

//BADD_653 replaced by BADD_1157

//BADD_652 replaced by BADD_1156

//BADD_651 replaced by BADD_1155

//BADD_650 replaced by BADD_1154

//BADD_649 replaced by BADD_1153

//BADD_648 replaced by BADD_1152

//BADD_647 replaced by BADD_1151

//BADD_646 replaced by BADD_1150

//BADD_645 replaced by BADD_1149

//BADD_644 replaced by BADD_1148

//BADD_643 replaced by BADD_1147

//BADD_642 replaced by BADD_1146

//BADD_641 replaced by BADD_1145

//BADD_640 replaced by BADD_1144

//BADD_639 replaced by BADD_1143

//BADD_638 replaced by BADD_1142

//BADD_637 replaced by BADD_1141

//BADD_636 replaced by BADD_1140

//BADD_635 replaced by BADD_1139

//BADD_634 replaced by BADD_1138

//BADD_633 replaced by BADD_1137

//BADD_632 replaced by BADD_1136

//BADD_631 replaced by BADD_1135

//BADD_630 replaced by BADD_1134

//BADD_629 replaced by BADD_1133

//BADD_628 replaced by BADD_1132

//BADD_627 replaced by BADD_1131

//BADD_626 replaced by BADD_1130

//BADD_625 replaced by BADD_1129

//BADD_624 replaced by BADD_1128

//BADD_623 replaced by BADD_1127

//BADD_622 replaced by BADD_1126

//BADD_621 replaced by BADD_1125

//KaratsubaCore_18 replaced by KaratsubaCore_35

//KaratsubaCore_19 replaced by KaratsubaCore_35

//FineReduction_46 replaced by FineReduction_53

//BADD_683 replaced by BADD_1124

//ADD_179 replaced by ADD_4223

//ADD_178 replaced by ADD_5756

//ADD_177 replaced by ADD_5756

//ADD_176 replaced by ADD_5756

//ADD_175 replaced by ADD_5756

//ADD_174 replaced by ADD_5756

//BADD_745 replaced by BADD_1186

//BADD_744 replaced by BADD_1185

//BADD_743 replaced by BADD_1184

//BADD_742 replaced by BADD_1183

//BADD_741 replaced by BADD_1182

//BADD_740 replaced by BADD_1181

//BADD_739 replaced by BADD_1180

//BADD_738 replaced by BADD_1179

//BADD_737 replaced by BADD_1178

//BADD_736 replaced by BADD_1177

//BADD_735 replaced by BADD_1176

//BADD_734 replaced by BADD_1175

//BADD_733 replaced by BADD_1174

//BADD_732 replaced by BADD_1173

//BADD_731 replaced by BADD_1172

//BADD_730 replaced by BADD_1171

//BADD_729 replaced by BADD_1170

//BADD_728 replaced by BADD_1169

//BADD_727 replaced by BADD_1168

//BADD_726 replaced by BADD_1167

//BADD_725 replaced by BADD_1166

//BADD_724 replaced by BADD_1165

//BADD_723 replaced by BADD_1164

//BADD_722 replaced by BADD_1163

//BADD_721 replaced by BADD_1162

//BADD_720 replaced by BADD_1161

//BADD_719 replaced by BADD_1160

//BADD_718 replaced by BADD_1159

//BADD_717 replaced by BADD_1158

//BADD_716 replaced by BADD_1157

//BADD_715 replaced by BADD_1156

//BADD_714 replaced by BADD_1155

//BADD_713 replaced by BADD_1154

//BADD_712 replaced by BADD_1153

//BADD_711 replaced by BADD_1152

//BADD_710 replaced by BADD_1151

//BADD_709 replaced by BADD_1150

//BADD_708 replaced by BADD_1149

//BADD_707 replaced by BADD_1148

//BADD_706 replaced by BADD_1147

//BADD_705 replaced by BADD_1146

//BADD_704 replaced by BADD_1145

//BADD_703 replaced by BADD_1144

//BADD_702 replaced by BADD_1143

//BADD_701 replaced by BADD_1142

//BADD_700 replaced by BADD_1141

//BADD_699 replaced by BADD_1140

//BADD_698 replaced by BADD_1139

//BADD_697 replaced by BADD_1138

//BADD_696 replaced by BADD_1137

//BADD_695 replaced by BADD_1136

//BADD_694 replaced by BADD_1135

//BADD_693 replaced by BADD_1134

//BADD_692 replaced by BADD_1133

//BADD_691 replaced by BADD_1132

//BADD_690 replaced by BADD_1131

//BADD_689 replaced by BADD_1130

//BADD_688 replaced by BADD_1129

//BADD_687 replaced by BADD_1128

//BADD_686 replaced by BADD_1127

//BADD_685 replaced by BADD_1126

//BADD_684 replaced by BADD_1125

//KaratsubaCore_20 replaced by KaratsubaCore_35

//KaratsubaCore_21 replaced by KaratsubaCore_35

//FineReduction_47 replaced by FineReduction_53

//BADD_746 replaced by BADD_1124

//ADD_185 replaced by ADD_4223

//ADD_184 replaced by ADD_5756

//ADD_183 replaced by ADD_5756

//ADD_182 replaced by ADD_5756

//ADD_181 replaced by ADD_5756

//ADD_180 replaced by ADD_5756

//BADD_808 replaced by BADD_1186

//BADD_807 replaced by BADD_1185

//BADD_806 replaced by BADD_1184

//BADD_805 replaced by BADD_1183

//BADD_804 replaced by BADD_1182

//BADD_803 replaced by BADD_1181

//BADD_802 replaced by BADD_1180

//BADD_801 replaced by BADD_1179

//BADD_800 replaced by BADD_1178

//BADD_799 replaced by BADD_1177

//BADD_798 replaced by BADD_1176

//BADD_797 replaced by BADD_1175

//BADD_796 replaced by BADD_1174

//BADD_795 replaced by BADD_1173

//BADD_794 replaced by BADD_1172

//BADD_793 replaced by BADD_1171

//BADD_792 replaced by BADD_1170

//BADD_791 replaced by BADD_1169

//BADD_790 replaced by BADD_1168

//BADD_789 replaced by BADD_1167

//BADD_788 replaced by BADD_1166

//BADD_787 replaced by BADD_1165

//BADD_786 replaced by BADD_1164

//BADD_785 replaced by BADD_1163

//BADD_784 replaced by BADD_1162

//BADD_783 replaced by BADD_1161

//BADD_782 replaced by BADD_1160

//BADD_781 replaced by BADD_1159

//BADD_780 replaced by BADD_1158

//BADD_779 replaced by BADD_1157

//BADD_778 replaced by BADD_1156

//BADD_777 replaced by BADD_1155

//BADD_776 replaced by BADD_1154

//BADD_775 replaced by BADD_1153

//BADD_774 replaced by BADD_1152

//BADD_773 replaced by BADD_1151

//BADD_772 replaced by BADD_1150

//BADD_771 replaced by BADD_1149

//BADD_770 replaced by BADD_1148

//BADD_769 replaced by BADD_1147

//BADD_768 replaced by BADD_1146

//BADD_767 replaced by BADD_1145

//BADD_766 replaced by BADD_1144

//BADD_765 replaced by BADD_1143

//BADD_764 replaced by BADD_1142

//BADD_763 replaced by BADD_1141

//BADD_762 replaced by BADD_1140

//BADD_761 replaced by BADD_1139

//BADD_760 replaced by BADD_1138

//BADD_759 replaced by BADD_1137

//BADD_758 replaced by BADD_1136

//BADD_757 replaced by BADD_1135

//BADD_756 replaced by BADD_1134

//BADD_755 replaced by BADD_1133

//BADD_754 replaced by BADD_1132

//BADD_753 replaced by BADD_1131

//BADD_752 replaced by BADD_1130

//BADD_751 replaced by BADD_1129

//BADD_750 replaced by BADD_1128

//BADD_749 replaced by BADD_1127

//BADD_748 replaced by BADD_1126

//BADD_747 replaced by BADD_1125

//KaratsubaCore_22 replaced by KaratsubaCore_35

//KaratsubaCore_23 replaced by KaratsubaCore_35

//FineReduction_48 replaced by FineReduction_53

//BADD_809 replaced by BADD_1124

//ADD_191 replaced by ADD_4223

//ADD_190 replaced by ADD_5756

//ADD_189 replaced by ADD_5756

//ADD_188 replaced by ADD_5756

//ADD_187 replaced by ADD_5756

//ADD_186 replaced by ADD_5756

//BADD_871 replaced by BADD_1186

//BADD_870 replaced by BADD_1185

//BADD_869 replaced by BADD_1184

//BADD_868 replaced by BADD_1183

//BADD_867 replaced by BADD_1182

//BADD_866 replaced by BADD_1181

//BADD_865 replaced by BADD_1180

//BADD_864 replaced by BADD_1179

//BADD_863 replaced by BADD_1178

//BADD_862 replaced by BADD_1177

//BADD_861 replaced by BADD_1176

//BADD_860 replaced by BADD_1175

//BADD_859 replaced by BADD_1174

//BADD_858 replaced by BADD_1173

//BADD_857 replaced by BADD_1172

//BADD_856 replaced by BADD_1171

//BADD_855 replaced by BADD_1170

//BADD_854 replaced by BADD_1169

//BADD_853 replaced by BADD_1168

//BADD_852 replaced by BADD_1167

//BADD_851 replaced by BADD_1166

//BADD_850 replaced by BADD_1165

//BADD_849 replaced by BADD_1164

//BADD_848 replaced by BADD_1163

//BADD_847 replaced by BADD_1162

//BADD_846 replaced by BADD_1161

//BADD_845 replaced by BADD_1160

//BADD_844 replaced by BADD_1159

//BADD_843 replaced by BADD_1158

//BADD_842 replaced by BADD_1157

//BADD_841 replaced by BADD_1156

//BADD_840 replaced by BADD_1155

//BADD_839 replaced by BADD_1154

//BADD_838 replaced by BADD_1153

//BADD_837 replaced by BADD_1152

//BADD_836 replaced by BADD_1151

//BADD_835 replaced by BADD_1150

//BADD_834 replaced by BADD_1149

//BADD_833 replaced by BADD_1148

//BADD_832 replaced by BADD_1147

//BADD_831 replaced by BADD_1146

//BADD_830 replaced by BADD_1145

//BADD_829 replaced by BADD_1144

//BADD_828 replaced by BADD_1143

//BADD_827 replaced by BADD_1142

//BADD_826 replaced by BADD_1141

//BADD_825 replaced by BADD_1140

//BADD_824 replaced by BADD_1139

//BADD_823 replaced by BADD_1138

//BADD_822 replaced by BADD_1137

//BADD_821 replaced by BADD_1136

//BADD_820 replaced by BADD_1135

//BADD_819 replaced by BADD_1134

//BADD_818 replaced by BADD_1133

//BADD_817 replaced by BADD_1132

//BADD_816 replaced by BADD_1131

//BADD_815 replaced by BADD_1130

//BADD_814 replaced by BADD_1129

//BADD_813 replaced by BADD_1128

//BADD_812 replaced by BADD_1127

//BADD_811 replaced by BADD_1126

//BADD_810 replaced by BADD_1125

//KaratsubaCore_24 replaced by KaratsubaCore_35

//KaratsubaCore_25 replaced by KaratsubaCore_35

//FineReduction_49 replaced by FineReduction_53

//BADD_872 replaced by BADD_1124

//ADD_197 replaced by ADD_4223

//ADD_196 replaced by ADD_5756

//ADD_195 replaced by ADD_5756

//ADD_194 replaced by ADD_5756

//ADD_193 replaced by ADD_5756

//ADD_192 replaced by ADD_5756

//BADD_934 replaced by BADD_1186

//BADD_933 replaced by BADD_1185

//BADD_932 replaced by BADD_1184

//BADD_931 replaced by BADD_1183

//BADD_930 replaced by BADD_1182

//BADD_929 replaced by BADD_1181

//BADD_928 replaced by BADD_1180

//BADD_927 replaced by BADD_1179

//BADD_926 replaced by BADD_1178

//BADD_925 replaced by BADD_1177

//BADD_924 replaced by BADD_1176

//BADD_923 replaced by BADD_1175

//BADD_922 replaced by BADD_1174

//BADD_921 replaced by BADD_1173

//BADD_920 replaced by BADD_1172

//BADD_919 replaced by BADD_1171

//BADD_918 replaced by BADD_1170

//BADD_917 replaced by BADD_1169

//BADD_916 replaced by BADD_1168

//BADD_915 replaced by BADD_1167

//BADD_914 replaced by BADD_1166

//BADD_913 replaced by BADD_1165

//BADD_912 replaced by BADD_1164

//BADD_911 replaced by BADD_1163

//BADD_910 replaced by BADD_1162

//BADD_909 replaced by BADD_1161

//BADD_908 replaced by BADD_1160

//BADD_907 replaced by BADD_1159

//BADD_906 replaced by BADD_1158

//BADD_905 replaced by BADD_1157

//BADD_904 replaced by BADD_1156

//BADD_903 replaced by BADD_1155

//BADD_902 replaced by BADD_1154

//BADD_901 replaced by BADD_1153

//BADD_900 replaced by BADD_1152

//BADD_899 replaced by BADD_1151

//BADD_898 replaced by BADD_1150

//BADD_897 replaced by BADD_1149

//BADD_896 replaced by BADD_1148

//BADD_895 replaced by BADD_1147

//BADD_894 replaced by BADD_1146

//BADD_893 replaced by BADD_1145

//BADD_892 replaced by BADD_1144

//BADD_891 replaced by BADD_1143

//BADD_890 replaced by BADD_1142

//BADD_889 replaced by BADD_1141

//BADD_888 replaced by BADD_1140

//BADD_887 replaced by BADD_1139

//BADD_886 replaced by BADD_1138

//BADD_885 replaced by BADD_1137

//BADD_884 replaced by BADD_1136

//BADD_883 replaced by BADD_1135

//BADD_882 replaced by BADD_1134

//BADD_881 replaced by BADD_1133

//BADD_880 replaced by BADD_1132

//BADD_879 replaced by BADD_1131

//BADD_878 replaced by BADD_1130

//BADD_877 replaced by BADD_1129

//BADD_876 replaced by BADD_1128

//BADD_875 replaced by BADD_1127

//BADD_874 replaced by BADD_1126

//BADD_873 replaced by BADD_1125

//KaratsubaCore_26 replaced by KaratsubaCore_35

//KaratsubaCore_27 replaced by KaratsubaCore_35

//FineReduction_50 replaced by FineReduction_53

//BADD_935 replaced by BADD_1124

//ADD_203 replaced by ADD_4223

//ADD_202 replaced by ADD_5756

//ADD_201 replaced by ADD_5756

//ADD_200 replaced by ADD_5756

//ADD_199 replaced by ADD_5756

//ADD_198 replaced by ADD_5756

//BADD_997 replaced by BADD_1186

//BADD_996 replaced by BADD_1185

//BADD_995 replaced by BADD_1184

//BADD_994 replaced by BADD_1183

//BADD_993 replaced by BADD_1182

//BADD_992 replaced by BADD_1181

//BADD_991 replaced by BADD_1180

//BADD_990 replaced by BADD_1179

//BADD_989 replaced by BADD_1178

//BADD_988 replaced by BADD_1177

//BADD_987 replaced by BADD_1176

//BADD_986 replaced by BADD_1175

//BADD_985 replaced by BADD_1174

//BADD_984 replaced by BADD_1173

//BADD_983 replaced by BADD_1172

//BADD_982 replaced by BADD_1171

//BADD_981 replaced by BADD_1170

//BADD_980 replaced by BADD_1169

//BADD_979 replaced by BADD_1168

//BADD_978 replaced by BADD_1167

//BADD_977 replaced by BADD_1166

//BADD_976 replaced by BADD_1165

//BADD_975 replaced by BADD_1164

//BADD_974 replaced by BADD_1163

//BADD_973 replaced by BADD_1162

//BADD_972 replaced by BADD_1161

//BADD_971 replaced by BADD_1160

//BADD_970 replaced by BADD_1159

//BADD_969 replaced by BADD_1158

//BADD_968 replaced by BADD_1157

//BADD_967 replaced by BADD_1156

//BADD_966 replaced by BADD_1155

//BADD_965 replaced by BADD_1154

//BADD_964 replaced by BADD_1153

//BADD_963 replaced by BADD_1152

//BADD_962 replaced by BADD_1151

//BADD_961 replaced by BADD_1150

//BADD_960 replaced by BADD_1149

//BADD_959 replaced by BADD_1148

//BADD_958 replaced by BADD_1147

//BADD_957 replaced by BADD_1146

//BADD_956 replaced by BADD_1145

//BADD_955 replaced by BADD_1144

//BADD_954 replaced by BADD_1143

//BADD_953 replaced by BADD_1142

//BADD_952 replaced by BADD_1141

//BADD_951 replaced by BADD_1140

//BADD_950 replaced by BADD_1139

//BADD_949 replaced by BADD_1138

//BADD_948 replaced by BADD_1137

//BADD_947 replaced by BADD_1136

//BADD_946 replaced by BADD_1135

//BADD_945 replaced by BADD_1134

//BADD_944 replaced by BADD_1133

//BADD_943 replaced by BADD_1132

//BADD_942 replaced by BADD_1131

//BADD_941 replaced by BADD_1130

//BADD_940 replaced by BADD_1129

//BADD_939 replaced by BADD_1128

//BADD_938 replaced by BADD_1127

//BADD_937 replaced by BADD_1126

//BADD_936 replaced by BADD_1125

//KaratsubaCore_28 replaced by KaratsubaCore_35

//KaratsubaCore_29 replaced by KaratsubaCore_35

//FineReduction_51 replaced by FineReduction_53

//BADD_998 replaced by BADD_1124

//ADD_209 replaced by ADD_4223

//ADD_208 replaced by ADD_5756

//ADD_207 replaced by ADD_5756

//ADD_206 replaced by ADD_5756

//ADD_205 replaced by ADD_5756

//ADD_204 replaced by ADD_5756

//BADD_1060 replaced by BADD_1186

//BADD_1059 replaced by BADD_1185

//BADD_1058 replaced by BADD_1184

//BADD_1057 replaced by BADD_1183

//BADD_1056 replaced by BADD_1182

//BADD_1055 replaced by BADD_1181

//BADD_1054 replaced by BADD_1180

//BADD_1053 replaced by BADD_1179

//BADD_1052 replaced by BADD_1178

//BADD_1051 replaced by BADD_1177

//BADD_1050 replaced by BADD_1176

//BADD_1049 replaced by BADD_1175

//BADD_1048 replaced by BADD_1174

//BADD_1047 replaced by BADD_1173

//BADD_1046 replaced by BADD_1172

//BADD_1045 replaced by BADD_1171

//BADD_1044 replaced by BADD_1170

//BADD_1043 replaced by BADD_1169

//BADD_1042 replaced by BADD_1168

//BADD_1041 replaced by BADD_1167

//BADD_1040 replaced by BADD_1166

//BADD_1039 replaced by BADD_1165

//BADD_1038 replaced by BADD_1164

//BADD_1037 replaced by BADD_1163

//BADD_1036 replaced by BADD_1162

//BADD_1035 replaced by BADD_1161

//BADD_1034 replaced by BADD_1160

//BADD_1033 replaced by BADD_1159

//BADD_1032 replaced by BADD_1158

//BADD_1031 replaced by BADD_1157

//BADD_1030 replaced by BADD_1156

//BADD_1029 replaced by BADD_1155

//BADD_1028 replaced by BADD_1154

//BADD_1027 replaced by BADD_1153

//BADD_1026 replaced by BADD_1152

//BADD_1025 replaced by BADD_1151

//BADD_1024 replaced by BADD_1150

//BADD_1023 replaced by BADD_1149

//BADD_1022 replaced by BADD_1148

//BADD_1021 replaced by BADD_1147

//BADD_1020 replaced by BADD_1146

//BADD_1019 replaced by BADD_1145

//BADD_1018 replaced by BADD_1144

//BADD_1017 replaced by BADD_1143

//BADD_1016 replaced by BADD_1142

//BADD_1015 replaced by BADD_1141

//BADD_1014 replaced by BADD_1140

//BADD_1013 replaced by BADD_1139

//BADD_1012 replaced by BADD_1138

//BADD_1011 replaced by BADD_1137

//BADD_1010 replaced by BADD_1136

//BADD_1009 replaced by BADD_1135

//BADD_1008 replaced by BADD_1134

//BADD_1007 replaced by BADD_1133

//BADD_1006 replaced by BADD_1132

//BADD_1005 replaced by BADD_1131

//BADD_1004 replaced by BADD_1130

//BADD_1003 replaced by BADD_1129

//BADD_1002 replaced by BADD_1128

//BADD_1001 replaced by BADD_1127

//BADD_1000 replaced by BADD_1126

//BADD_999 replaced by BADD_1125

//KaratsubaCore_30 replaced by KaratsubaCore_35

//KaratsubaCore_31 replaced by KaratsubaCore_35

//FineReduction_52 replaced by FineReduction_53

//BADD_1061 replaced by BADD_1124

//ADD_215 replaced by ADD_4223

//ADD_214 replaced by ADD_5756

//ADD_213 replaced by ADD_5756

//ADD_212 replaced by ADD_5756

//ADD_211 replaced by ADD_5756

//ADD_210 replaced by ADD_5756

//BADD_1123 replaced by BADD_1186

//BADD_1122 replaced by BADD_1185

//BADD_1121 replaced by BADD_1184

//BADD_1120 replaced by BADD_1183

//BADD_1119 replaced by BADD_1182

//BADD_1118 replaced by BADD_1181

//BADD_1117 replaced by BADD_1180

//BADD_1116 replaced by BADD_1179

//BADD_1115 replaced by BADD_1178

//BADD_1114 replaced by BADD_1177

//BADD_1113 replaced by BADD_1176

//BADD_1112 replaced by BADD_1175

//BADD_1111 replaced by BADD_1174

//BADD_1110 replaced by BADD_1173

//BADD_1109 replaced by BADD_1172

//BADD_1108 replaced by BADD_1171

//BADD_1107 replaced by BADD_1170

//BADD_1106 replaced by BADD_1169

//BADD_1105 replaced by BADD_1168

//BADD_1104 replaced by BADD_1167

//BADD_1103 replaced by BADD_1166

//BADD_1102 replaced by BADD_1165

//BADD_1101 replaced by BADD_1164

//BADD_1100 replaced by BADD_1163

//BADD_1099 replaced by BADD_1162

//BADD_1098 replaced by BADD_1161

//BADD_1097 replaced by BADD_1160

//BADD_1096 replaced by BADD_1159

//BADD_1095 replaced by BADD_1158

//BADD_1094 replaced by BADD_1157

//BADD_1093 replaced by BADD_1156

//BADD_1092 replaced by BADD_1155

//BADD_1091 replaced by BADD_1154

//BADD_1090 replaced by BADD_1153

//BADD_1089 replaced by BADD_1152

//BADD_1088 replaced by BADD_1151

//BADD_1087 replaced by BADD_1150

//BADD_1086 replaced by BADD_1149

//BADD_1085 replaced by BADD_1148

//BADD_1084 replaced by BADD_1147

//BADD_1083 replaced by BADD_1146

//BADD_1082 replaced by BADD_1145

//BADD_1081 replaced by BADD_1144

//BADD_1080 replaced by BADD_1143

//BADD_1079 replaced by BADD_1142

//BADD_1078 replaced by BADD_1141

//BADD_1077 replaced by BADD_1140

//BADD_1076 replaced by BADD_1139

//BADD_1075 replaced by BADD_1138

//BADD_1074 replaced by BADD_1137

//BADD_1073 replaced by BADD_1136

//BADD_1072 replaced by BADD_1135

//BADD_1071 replaced by BADD_1134

//BADD_1070 replaced by BADD_1133

//BADD_1069 replaced by BADD_1132

//BADD_1068 replaced by BADD_1131

//BADD_1067 replaced by BADD_1130

//BADD_1066 replaced by BADD_1129

//BADD_1065 replaced by BADD_1128

//BADD_1064 replaced by BADD_1127

//BADD_1063 replaced by BADD_1126

//BADD_1062 replaced by BADD_1125

//KaratsubaCore_32 replaced by KaratsubaCore_35

//KaratsubaCore_33 replaced by KaratsubaCore_35

module FineReduction_53 (
  input      [377:0]  io_a,
  output     [376:0]  io_r,
  input               clk,
  input               resetn
);

  wire       [378:0]  singleAdd_add_io_s;
  wire       [376:0]  _zz__zz_io_r;
  wire       [376:0]  _zz__zz_io_r_1;
  reg        [63:0]   _zz_singleAdd_a;
  reg        [63:0]   _zz_singleAdd_a_1;
  reg        [63:0]   _zz_singleAdd_a_2;
  reg        [63:0]   _zz_singleAdd_a_3;
  reg        [63:0]   _zz_singleAdd_a_4;
  reg        [63:0]   _zz_singleAdd_a_5;
  reg        [63:0]   _zz_singleAdd_a_6;
  reg        [63:0]   _zz_singleAdd_a_7;
  reg        [63:0]   _zz_singleAdd_a_8;
  reg        [63:0]   _zz_singleAdd_a_9;
  reg        [63:0]   _zz_singleAdd_a_10;
  reg        [63:0]   _zz_singleAdd_a_11;
  reg        [63:0]   _zz_singleAdd_a_12;
  reg        [63:0]   _zz_singleAdd_a_13;
  reg        [63:0]   _zz_singleAdd_a_14;
  reg        [63:0]   _zz_singleAdd_a_15;
  reg        [63:0]   _zz_singleAdd_a_16;
  reg        [63:0]   _zz_singleAdd_a_17;
  reg        [63:0]   _zz_singleAdd_a_18;
  reg        [63:0]   _zz_singleAdd_a_19;
  reg        [57:0]   _zz_singleAdd_a_20;
  wire       [377:0]  singleAdd_a;
  reg        [376:0]  _zz_io_r;

  assign _zz__zz_io_r = singleAdd_add_io_s[376:0];
  assign _zz__zz_io_r_1 = singleAdd_a[376:0];
  BADD_1306 singleAdd_add (
    .io_a   (io_a[377:0]                                                                                         ), //i
    .io_b   (378'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001), //i
    .io_c   (1'b0                                                                                                ), //i
    .io_s   (singleAdd_add_io_s[378:0]                                                                           ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  assign singleAdd_a = {_zz_singleAdd_a_20,{_zz_singleAdd_a_19,{_zz_singleAdd_a_17,{_zz_singleAdd_a_14,{_zz_singleAdd_a_10,_zz_singleAdd_a_5}}}}};
  assign io_r = _zz_io_r;
  always @(posedge clk) begin
    _zz_singleAdd_a <= io_a[63 : 0];
    _zz_singleAdd_a_1 <= _zz_singleAdd_a;
    _zz_singleAdd_a_2 <= _zz_singleAdd_a_1;
    _zz_singleAdd_a_3 <= _zz_singleAdd_a_2;
    _zz_singleAdd_a_4 <= _zz_singleAdd_a_3;
    _zz_singleAdd_a_5 <= _zz_singleAdd_a_4;
    _zz_singleAdd_a_6 <= io_a[127 : 64];
    _zz_singleAdd_a_7 <= _zz_singleAdd_a_6;
    _zz_singleAdd_a_8 <= _zz_singleAdd_a_7;
    _zz_singleAdd_a_9 <= _zz_singleAdd_a_8;
    _zz_singleAdd_a_10 <= _zz_singleAdd_a_9;
    _zz_singleAdd_a_11 <= io_a[191 : 128];
    _zz_singleAdd_a_12 <= _zz_singleAdd_a_11;
    _zz_singleAdd_a_13 <= _zz_singleAdd_a_12;
    _zz_singleAdd_a_14 <= _zz_singleAdd_a_13;
    _zz_singleAdd_a_15 <= io_a[255 : 192];
    _zz_singleAdd_a_16 <= _zz_singleAdd_a_15;
    _zz_singleAdd_a_17 <= _zz_singleAdd_a_16;
    _zz_singleAdd_a_18 <= io_a[319 : 256];
    _zz_singleAdd_a_19 <= _zz_singleAdd_a_18;
    _zz_singleAdd_a_20 <= io_a[377 : 320];
    _zz_io_r <= (singleAdd_a[377] ? _zz__zz_io_r : _zz__zz_io_r_1);
  end


endmodule

module BADD_1124 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  input               io_c,
  output     [378:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [57:0]   adder_adds_5_io_A_0;
  wire       [57:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [58:0]   adder_adds_5_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [63:0]   _zz_io_A_0_6;
  reg        [63:0]   _zz_io_A_0_7;
  reg        [63:0]   _zz_io_A_0_8;
  reg        [63:0]   _zz_io_A_0_9;
  reg        [57:0]   _zz_io_A_0_10;
  reg        [57:0]   _zz_io_A_0_11;
  reg        [57:0]   _zz_io_A_0_12;
  reg        [57:0]   _zz_io_A_0_13;
  reg        [57:0]   _zz_io_A_0_14;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [63:0]   _zz_io_A_1_6;
  reg        [63:0]   _zz_io_A_1_7;
  reg        [63:0]   _zz_io_A_1_8;
  reg        [63:0]   _zz_io_A_1_9;
  reg        [57:0]   _zz_io_A_1_10;
  reg        [57:0]   _zz_io_A_1_11;
  reg        [57:0]   _zz_io_A_1_12;
  reg        [57:0]   _zz_io_A_1_13;
  reg        [57:0]   _zz_io_A_1_14;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [57:0]   _zz_io_s_6;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_5761 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[57:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[57:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[58:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_5_io_A_0 = _zz_io_A_0_14;
  assign adder_adds_0_io_A_1 = (~ io_b[63 : 0]);
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign adder_adds_5_io_A_1 = _zz_io_A_1_14;
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[319 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_0_10 <= io_a[377 : 320];
    _zz_io_A_0_11 <= _zz_io_A_0_10;
    _zz_io_A_0_12 <= _zz_io_A_0_11;
    _zz_io_A_0_13 <= _zz_io_A_0_12;
    _zz_io_A_0_14 <= _zz_io_A_0_13;
    _zz_io_A_1 <= (~ io_b[127 : 64]);
    _zz_io_A_1_1 <= (~ io_b[191 : 128]);
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= (~ io_b[255 : 192]);
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= (~ io_b[319 : 256]);
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_A_1_10 <= (~ io_b[377 : 320]);
    _zz_io_A_1_11 <= _zz_io_A_1_10;
    _zz_io_A_1_12 <= _zz_io_A_1_11;
    _zz_io_A_1_13 <= _zz_io_A_1_12;
    _zz_io_A_1_14 <= _zz_io_A_1_13;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= (! adder_adds_5_io_S[58]);
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[57 : 0];
  end


endmodule

//ADD_221 replaced by ADD_4223

//ADD_220 replaced by ADD_5756

//ADD_219 replaced by ADD_5756

//ADD_218 replaced by ADD_5756

//ADD_217 replaced by ADD_5756

//ADD_216 replaced by ADD_5756

module BADD_1186 (
  input      [378:0]  io_a,
  input      [378:0]  io_b,
  input               io_c,
  output     [379:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [58:0]   adder_adds_5_io_A_0;
  wire       [58:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [59:0]   adder_adds_5_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  reg        [58:0]   _zz_io_s_21;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = io_a[127 : 64];
  assign adder_adds_2_io_A_0 = io_a[191 : 128];
  assign adder_adds_3_io_A_0 = io_a[255 : 192];
  assign adder_adds_4_io_A_0 = io_a[319 : 256];
  assign adder_adds_5_io_A_0 = io_a[378 : 320];
  assign adder_adds_0_io_A_1 = (~ io_b[63 : 0]);
  assign adder_adds_1_io_A_1 = (~ io_b[127 : 64]);
  assign adder_adds_2_io_A_1 = (~ io_b[191 : 128]);
  assign adder_adds_3_io_A_1 = (~ io_b[255 : 192]);
  assign adder_adds_4_io_A_1 = (~ io_b[319 : 256]);
  assign adder_adds_5_io_A_1 = (~ io_b[378 : 320]);
  assign io_s = {_zz_io_s,{_zz_io_s_21,{_zz_io_s_20,{_zz_io_s_18,{_zz_io_s_15,{_zz_io_s_11,_zz_io_s_6}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= (! adder_adds_5_io_S[59]);
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_8 <= _zz_io_s_7;
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_21 <= adder_adds_5_io_S[58 : 0];
  end


endmodule

module BADD_1185 (
  input      [120:0]  io_a,
  input      [120:0]  io_b,
  input               io_c,
  output     [121:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [61:0]   adder_adds_0_io_A_0;
  wire       [61:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [62:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [61:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4226 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[61:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[61:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[62:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[61 : 0];
  assign adder_adds_1_io_A_0 = io_a[120 : 62];
  assign adder_adds_0_io_A_1 = io_b[61 : 0];
  assign adder_adds_1_io_A_1 = io_b[120 : 62];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[62];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[61 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1184 (
  input      [36:0]   io_a,
  input      [36:0]   io_b,
  input               io_c,
  output     [37:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [36:0]   adder_adds_0_io_A_0;
  wire       [36:0]   adder_adds_0_io_A_1;
  wire       [37:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [36:0]   _zz_io_s_1;

  ADD_4055 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[36:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[36:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[37:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[36 : 0];
  assign adder_adds_0_io_A_1 = io_b[36 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[37];
    _zz_io_s_1 <= adder_adds_0_io_S[36 : 0];
  end


endmodule

module BADD_1183 (
  input      [9:0]    io_a,
  input      [9:0]    io_b,
  input               io_c,
  output     [10:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [9:0]    adder_adds_0_io_A_0;
  wire       [9:0]    adder_adds_0_io_A_1;
  wire       [10:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [9:0]    _zz_io_s_1;

  ADD_4057 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[9:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[9:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[10:0] )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[9 : 0];
  assign adder_adds_0_io_A_1 = io_b[9 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[10];
    _zz_io_s_1 <= adder_adds_0_io_S[9 : 0];
  end


endmodule

module BADD_1182 (
  input      [68:0]   io_a,
  input      [68:0]   io_b,
  input               io_c,
  output     [69:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [9:0]    adder_adds_0_io_A_0;
  wire       [9:0]    adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [10:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [9:0]    _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4057 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[9:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[9:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[10:0] )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[9 : 0];
  assign adder_adds_1_io_A_0 = io_a[68 : 10];
  assign adder_adds_0_io_A_1 = io_b[9 : 0];
  assign adder_adds_1_io_A_1 = io_b[68 : 10];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[10];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[9 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1181 (
  input      [58:0]   io_a,
  input      [58:0]   io_b,
  input               io_c,
  output     [59:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [58:0]   adder_adds_0_io_A_0;
  wire       [58:0]   adder_adds_0_io_A_1;
  wire       [59:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [58:0]   _zz_io_s_1;

  ADD_4223 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[58:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[58 : 0];
  assign adder_adds_0_io_A_1 = io_b[58 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[58 : 0];
  end


endmodule

module BADD_1180 (
  input      [54:0]   io_a,
  input      [54:0]   io_b,
  input               io_c,
  output     [55:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [54:0]   adder_adds_0_io_A_0;
  wire       [54:0]   adder_adds_0_io_A_1;
  wire       [55:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [54:0]   _zz_io_s_1;

  ADD_4060 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[54:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[54:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[55:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[54 : 0];
  assign adder_adds_0_io_A_1 = io_b[54 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[55];
    _zz_io_s_1 <= adder_adds_0_io_S[54 : 0];
  end


endmodule

module BADD_1179 (
  input      [63:0]   io_a,
  input      [63:0]   io_b,
  input               io_c,
  output     [64:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [4:0]    adder_adds_0_io_A_0;
  wire       [4:0]    adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [5:0]    adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [4:0]    _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_11560 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[4:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[4:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[5:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[4 : 0];
  assign adder_adds_1_io_A_0 = io_a[63 : 5];
  assign adder_adds_0_io_A_1 = io_b[4 : 0];
  assign adder_adds_1_io_A_1 = io_b[63 : 5];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[5];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[4 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1178 (
  input      [84:0]   io_a,
  input      [84:0]   io_b,
  input               io_c,
  output     [85:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [25:0]   adder_adds_0_io_A_0;
  wire       [25:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [26:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [25:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4196 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[25:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[25:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[26:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[25 : 0];
  assign adder_adds_1_io_A_0 = io_a[84 : 26];
  assign adder_adds_0_io_A_1 = io_b[25 : 0];
  assign adder_adds_1_io_A_1 = io_b[84 : 26];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[26];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[25 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1177 (
  input      [74:0]   io_a,
  input      [74:0]   io_b,
  input               io_c,
  output     [75:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [15:0]   adder_adds_0_io_A_0;
  wire       [15:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [16:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [15:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4132 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[15:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[15:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[16:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[15 : 0];
  assign adder_adds_1_io_A_0 = io_a[74 : 16];
  assign adder_adds_0_io_A_1 = io_b[15 : 0];
  assign adder_adds_1_io_A_1 = io_b[74 : 16];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[16];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[15 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1176 (
  input      [96:0]   io_a,
  input      [96:0]   io_b,
  input               io_c,
  output     [97:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [37:0]   adder_adds_0_io_A_0;
  wire       [37:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [38:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [37:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4067 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[37:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[37:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[38:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[37 : 0];
  assign adder_adds_1_io_A_0 = io_a[96 : 38];
  assign adder_adds_0_io_A_1 = io_b[37 : 0];
  assign adder_adds_1_io_A_1 = io_b[96 : 38];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[38];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[37 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1175 (
  input      [189:0]  io_a,
  input      [189:0]  io_b,
  input               io_c,
  output     [190:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [2:0]    adder_adds_0_io_A_0;
  wire       [2:0]    adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [3:0]    adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [2:0]    _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_11592 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[2:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[2:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[3:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[2 : 0];
  assign adder_adds_1_io_A_0 = io_a[66 : 3];
  assign adder_adds_2_io_A_0 = io_a[130 : 67];
  assign adder_adds_3_io_A_0 = io_a[189 : 131];
  assign adder_adds_0_io_A_1 = io_b[2 : 0];
  assign adder_adds_1_io_A_1 = io_b[66 : 3];
  assign adder_adds_2_io_A_1 = io_b[130 : 67];
  assign adder_adds_3_io_A_1 = io_b[189 : 131];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[3];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[2 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1174 (
  input      [145:0]  io_a,
  input      [145:0]  io_b,
  input               io_c,
  output     [146:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [22:0]   adder_adds_0_io_A_0;
  wire       [22:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [23:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [22:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4168 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[22:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[22:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[23:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[22 : 0];
  assign adder_adds_1_io_A_0 = io_a[86 : 23];
  assign adder_adds_2_io_A_0 = io_a[145 : 87];
  assign adder_adds_0_io_A_1 = io_b[22 : 0];
  assign adder_adds_1_io_A_1 = io_b[86 : 23];
  assign adder_adds_2_io_A_1 = io_b[145 : 87];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[23];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[22 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1173 (
  input      [129:0]  io_a,
  input      [129:0]  io_b,
  input               io_c,
  output     [130:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [6:0]    adder_adds_0_io_A_0;
  wire       [6:0]    adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [7:0]    adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [6:0]    _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4076 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[6:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[6:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[7:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[6 : 0];
  assign adder_adds_1_io_A_0 = io_a[70 : 7];
  assign adder_adds_2_io_A_0 = io_a[129 : 71];
  assign adder_adds_0_io_A_1 = io_b[6 : 0];
  assign adder_adds_1_io_A_1 = io_b[70 : 7];
  assign adder_adds_2_io_A_1 = io_b[129 : 71];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[7];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[6 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1172 (
  input      [125:0]  io_a,
  input      [125:0]  io_b,
  input               io_c,
  output     [126:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [2:0]    adder_adds_0_io_A_0;
  wire       [2:0]    adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [3:0]    adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [2:0]    _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_11592 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[2:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[2:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[3:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[2 : 0];
  assign adder_adds_1_io_A_0 = io_a[66 : 3];
  assign adder_adds_2_io_A_0 = io_a[125 : 67];
  assign adder_adds_0_io_A_1 = io_b[2 : 0];
  assign adder_adds_1_io_A_1 = io_b[66 : 3];
  assign adder_adds_2_io_A_1 = io_b[125 : 67];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[3];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[2 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1171 (
  input      [141:0]  io_a,
  input      [141:0]  io_b,
  input               io_c,
  output     [142:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [18:0]   adder_adds_0_io_A_0;
  wire       [18:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [19:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [18:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4106 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[18:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[18:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[19:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[18 : 0];
  assign adder_adds_1_io_A_0 = io_a[82 : 19];
  assign adder_adds_2_io_A_0 = io_a[141 : 83];
  assign adder_adds_0_io_A_1 = io_b[18 : 0];
  assign adder_adds_1_io_A_1 = io_b[82 : 19];
  assign adder_adds_2_io_A_1 = io_b[141 : 83];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[19];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[18 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1170 (
  input      [166:0]  io_a,
  input      [166:0]  io_b,
  input               io_c,
  output     [167:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [43:0]   adder_adds_0_io_A_0;
  wire       [43:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [44:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [43:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4085 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[43:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[43:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[44:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[43 : 0];
  assign adder_adds_1_io_A_0 = io_a[107 : 44];
  assign adder_adds_2_io_A_0 = io_a[166 : 108];
  assign adder_adds_0_io_A_1 = io_b[43 : 0];
  assign adder_adds_1_io_A_1 = io_b[107 : 44];
  assign adder_adds_2_io_A_1 = io_b[166 : 108];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[44];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[43 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1169 (
  input      [150:0]  io_a,
  input      [150:0]  io_b,
  input               io_c,
  output     [151:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [27:0]   adder_adds_0_io_A_0;
  wire       [27:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [28:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [27:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4158 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[27:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[27:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[28:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[27 : 0];
  assign adder_adds_1_io_A_0 = io_a[91 : 28];
  assign adder_adds_2_io_A_0 = io_a[150 : 92];
  assign adder_adds_0_io_A_1 = io_b[27 : 0];
  assign adder_adds_1_io_A_1 = io_b[91 : 28];
  assign adder_adds_2_io_A_1 = io_b[150 : 92];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[28];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[27 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1168 (
  input      [182:0]  io_a,
  input      [182:0]  io_b,
  input               io_c,
  output     [183:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [59:0]   adder_adds_0_io_A_0;
  wire       [59:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [60:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [59:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4091 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[59:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[59:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[60:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[59 : 0];
  assign adder_adds_1_io_A_0 = io_a[123 : 60];
  assign adder_adds_2_io_A_0 = io_a[182 : 124];
  assign adder_adds_0_io_A_1 = io_b[59 : 0];
  assign adder_adds_1_io_A_1 = io_b[123 : 60];
  assign adder_adds_2_io_A_1 = io_b[182 : 124];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[60];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[59 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1167 (
  input      [220:0]  io_a,
  input      [220:0]  io_b,
  input               io_c,
  output     [221:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [33:0]   adder_adds_0_io_A_0;
  wire       [33:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [34:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [33:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_4094 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[33:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[33:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[34:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[33 : 0];
  assign adder_adds_1_io_A_0 = io_a[97 : 34];
  assign adder_adds_2_io_A_0 = io_a[161 : 98];
  assign adder_adds_3_io_A_0 = io_a[220 : 162];
  assign adder_adds_0_io_A_1 = io_b[33 : 0];
  assign adder_adds_1_io_A_1 = io_b[97 : 34];
  assign adder_adds_2_io_A_1 = io_b[161 : 98];
  assign adder_adds_3_io_A_1 = io_b[220 : 162];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[34];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[33 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1166 (
  input      [200:0]  io_a,
  input      [200:0]  io_b,
  input               io_c,
  output     [201:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [13:0]   adder_adds_0_io_A_0;
  wire       [13:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [14:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [13:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_4145 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[13:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[13:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[14:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[13 : 0];
  assign adder_adds_1_io_A_0 = io_a[77 : 14];
  assign adder_adds_2_io_A_0 = io_a[141 : 78];
  assign adder_adds_3_io_A_0 = io_a[200 : 142];
  assign adder_adds_0_io_A_1 = io_b[13 : 0];
  assign adder_adds_1_io_A_1 = io_b[77 : 14];
  assign adder_adds_2_io_A_1 = io_b[141 : 78];
  assign adder_adds_3_io_A_1 = io_b[200 : 142];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[14];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[13 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1165 (
  input      [194:0]  io_a,
  input      [194:0]  io_b,
  input               io_c,
  output     [195:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [7:0]    adder_adds_0_io_A_0;
  wire       [7:0]    adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [8:0]    adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [7:0]    _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_4212 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[7:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[7:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[8:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[7 : 0];
  assign adder_adds_1_io_A_0 = io_a[71 : 8];
  assign adder_adds_2_io_A_0 = io_a[135 : 72];
  assign adder_adds_3_io_A_0 = io_a[194 : 136];
  assign adder_adds_0_io_A_1 = io_b[7 : 0];
  assign adder_adds_1_io_A_1 = io_b[71 : 8];
  assign adder_adds_2_io_A_1 = io_b[135 : 72];
  assign adder_adds_3_io_A_1 = io_b[194 : 136];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[8];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[7 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1164 (
  input      [205:0]  io_a,
  input      [205:0]  io_b,
  input               io_c,
  output     [206:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [18:0]   adder_adds_0_io_A_0;
  wire       [18:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [19:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [18:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_4106 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[18:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[18:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[19:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[18 : 0];
  assign adder_adds_1_io_A_0 = io_a[82 : 19];
  assign adder_adds_2_io_A_0 = io_a[146 : 83];
  assign adder_adds_3_io_A_0 = io_a[205 : 147];
  assign adder_adds_0_io_A_1 = io_b[18 : 0];
  assign adder_adds_1_io_A_1 = io_b[82 : 19];
  assign adder_adds_2_io_A_1 = io_b[146 : 83];
  assign adder_adds_3_io_A_1 = io_b[205 : 147];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[19];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[18 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1163 (
  input      [258:0]  io_a,
  input      [258:0]  io_b,
  input               io_c,
  output     [259:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [7:0]    adder_adds_0_io_A_0;
  wire       [7:0]    adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [58:0]   adder_adds_4_io_A_0;
  wire       [58:0]   adder_adds_4_io_A_1;
  wire       [8:0]    adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [59:0]   adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [7:0]    _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [58:0]   _zz_io_s_5;

  ADD_4212 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[7:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[7:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[8:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[7 : 0];
  assign adder_adds_1_io_A_0 = io_a[71 : 8];
  assign adder_adds_2_io_A_0 = io_a[135 : 72];
  assign adder_adds_3_io_A_0 = io_a[199 : 136];
  assign adder_adds_4_io_A_0 = io_a[258 : 200];
  assign adder_adds_0_io_A_1 = io_b[7 : 0];
  assign adder_adds_1_io_A_1 = io_b[71 : 8];
  assign adder_adds_2_io_A_1 = io_b[135 : 72];
  assign adder_adds_3_io_A_1 = io_b[199 : 136];
  assign adder_adds_4_io_A_1 = io_b[258 : 200];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[8];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_s <= adder_adds_4_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[7 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[58 : 0];
  end


endmodule

module BADD_1162 (
  input      [225:0]  io_a,
  input      [225:0]  io_b,
  input               io_c,
  output     [226:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [38:0]   adder_adds_0_io_A_0;
  wire       [38:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [39:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [38:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_4115 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[38:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[38:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[39:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[38 : 0];
  assign adder_adds_1_io_A_0 = io_a[102 : 39];
  assign adder_adds_2_io_A_0 = io_a[166 : 103];
  assign adder_adds_3_io_A_0 = io_a[225 : 167];
  assign adder_adds_0_io_A_1 = io_b[38 : 0];
  assign adder_adds_1_io_A_1 = io_b[102 : 39];
  assign adder_adds_2_io_A_1 = io_b[166 : 103];
  assign adder_adds_3_io_A_1 = io_b[225 : 167];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[39];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[38 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1161 (
  input      [267:0]  io_a,
  input      [267:0]  io_b,
  input               io_c,
  output     [268:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [16:0]   adder_adds_0_io_A_0;
  wire       [16:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [58:0]   adder_adds_4_io_A_0;
  wire       [58:0]   adder_adds_4_io_A_1;
  wire       [17:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [59:0]   adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [16:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [58:0]   _zz_io_s_5;

  ADD_4231 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[16:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[16:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[17:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[16 : 0];
  assign adder_adds_1_io_A_0 = io_a[80 : 17];
  assign adder_adds_2_io_A_0 = io_a[144 : 81];
  assign adder_adds_3_io_A_0 = io_a[208 : 145];
  assign adder_adds_4_io_A_0 = io_a[267 : 209];
  assign adder_adds_0_io_A_1 = io_b[16 : 0];
  assign adder_adds_1_io_A_1 = io_b[80 : 17];
  assign adder_adds_2_io_A_1 = io_b[144 : 81];
  assign adder_adds_3_io_A_1 = io_b[208 : 145];
  assign adder_adds_4_io_A_1 = io_b[267 : 209];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[17];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_s <= adder_adds_4_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[16 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[58 : 0];
  end


endmodule

module BADD_1160 (
  input      [4:0]    io_a,
  input      [4:0]    io_b,
  input               io_c,
  output     [5:0]    io_s,
  input               clk,
  input               resetn
);

  wire       [4:0]    adder_adds_0_io_A_0;
  wire       [4:0]    adder_adds_0_io_A_1;
  wire       [5:0]    adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [4:0]    _zz_io_s_1;

  ADD_11560 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[4:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[4:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[5:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[4 : 0];
  assign adder_adds_0_io_A_1 = io_b[4 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[5];
    _zz_io_s_1 <= adder_adds_0_io_S[4 : 0];
  end


endmodule

module BADD_1159 (
  input      [162:0]  io_a,
  input      [162:0]  io_b,
  input               io_c,
  output     [163:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [39:0]   adder_adds_0_io_A_0;
  wire       [39:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [40:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [39:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4125 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[39:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[39:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[40:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[39 : 0];
  assign adder_adds_1_io_A_0 = io_a[103 : 40];
  assign adder_adds_2_io_A_0 = io_a[162 : 104];
  assign adder_adds_0_io_A_1 = io_b[39 : 0];
  assign adder_adds_1_io_A_1 = io_b[103 : 40];
  assign adder_adds_2_io_A_1 = io_b[162 : 104];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[40];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[39 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1158 (
  input      [79:0]   io_a,
  input      [79:0]   io_b,
  input               io_c,
  output     [80:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [20:0]   adder_adds_0_io_A_0;
  wire       [20:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [21:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [20:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4131 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[20:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[20:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[21:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[20 : 0];
  assign adder_adds_1_io_A_0 = io_a[79 : 21];
  assign adder_adds_0_io_A_1 = io_b[20 : 0];
  assign adder_adds_1_io_A_1 = io_b[79 : 21];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[21];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[20 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1157 (
  input      [31:0]   io_a,
  input      [31:0]   io_b,
  input               io_c,
  output     [32:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [31:0]   adder_adds_0_io_A_0;
  wire       [31:0]   adder_adds_0_io_A_1;
  wire       [32:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [31:0]   _zz_io_s_1;

  ADD_4150 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[31:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[31:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[32:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[31 : 0];
  assign adder_adds_0_io_A_1 = io_b[31 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[32];
    _zz_io_s_1 <= adder_adds_0_io_S[31 : 0];
  end


endmodule

module BADD_1156 (
  input      [20:0]   io_a,
  input      [20:0]   io_b,
  input               io_c,
  output     [21:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [20:0]   adder_adds_0_io_A_0;
  wire       [20:0]   adder_adds_0_io_A_1;
  wire       [21:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [20:0]   _zz_io_s_1;

  ADD_4131 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[20:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[20:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[21:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[20 : 0];
  assign adder_adds_0_io_A_1 = io_b[20 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[21];
    _zz_io_s_1 <= adder_adds_0_io_S[20 : 0];
  end


endmodule

module BADD_1155 (
  input      [15:0]   io_a,
  input      [15:0]   io_b,
  input               io_c,
  output     [16:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [15:0]   adder_adds_0_io_A_0;
  wire       [15:0]   adder_adds_0_io_A_1;
  wire       [16:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [15:0]   _zz_io_s_1;

  ADD_4132 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[15:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[15:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[16:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[15 : 0];
  assign adder_adds_0_io_A_1 = io_b[15 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[16];
    _zz_io_s_1 <= adder_adds_0_io_S[15 : 0];
  end


endmodule

module BADD_1154 (
  input      [25:0]   io_a,
  input      [25:0]   io_b,
  input               io_c,
  output     [26:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [25:0]   adder_adds_0_io_A_0;
  wire       [25:0]   adder_adds_0_io_A_1;
  wire       [26:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [25:0]   _zz_io_s_1;

  ADD_4196 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[25:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[25:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[26:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[25 : 0];
  assign adder_adds_0_io_A_1 = io_b[25 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[26];
    _zz_io_s_1 <= adder_adds_0_io_S[25 : 0];
  end


endmodule

module BADD_1153 (
  input      [46:0]   io_a,
  input      [46:0]   io_b,
  input               io_c,
  output     [47:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [46:0]   adder_adds_0_io_A_0;
  wire       [46:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [46:0]   _zz_io_s_1;

  ADD_4134 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[46:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[46:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[47:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[46 : 0];
  assign adder_adds_0_io_A_1 = io_b[46 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[47];
    _zz_io_s_1 <= adder_adds_0_io_S[46 : 0];
  end


endmodule

module BADD_1152 (
  input      [42:0]   io_a,
  input      [42:0]   io_b,
  input               io_c,
  output     [43:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [42:0]   adder_adds_0_io_A_0;
  wire       [42:0]   adder_adds_0_io_A_1;
  wire       [43:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [42:0]   _zz_io_s_1;

  ADD_4139 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[42:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[42:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[43:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[42 : 0];
  assign adder_adds_0_io_A_1 = io_b[42 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[43];
    _zz_io_s_1 <= adder_adds_0_io_S[42 : 0];
  end


endmodule

module BADD_1151 (
  input      [50:0]   io_a,
  input      [50:0]   io_b,
  input               io_c,
  output     [51:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [50:0]   adder_adds_0_io_A_0;
  wire       [50:0]   adder_adds_0_io_A_1;
  wire       [51:0]   adder_adds_0_io_S;
  reg                 _zz_io_s;
  reg        [50:0]   _zz_io_s_1;

  ADD_4136 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[50:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[50:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[51:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[50 : 0];
  assign adder_adds_0_io_A_1 = io_b[50 : 0];
  assign io_s = {_zz_io_s,_zz_io_s_1};
  always @(posedge clk) begin
    _zz_io_s <= adder_adds_0_io_S[51];
    _zz_io_s_1 <= adder_adds_0_io_S[50 : 0];
  end


endmodule

module BADD_1150 (
  input      [111:0]  io_a,
  input      [111:0]  io_b,
  input               io_c,
  output     [112:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [52:0]   adder_adds_0_io_A_0;
  wire       [52:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [53:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [52:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4172 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[52:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[52:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[53:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[52 : 0];
  assign adder_adds_1_io_A_0 = io_a[111 : 53];
  assign adder_adds_0_io_A_1 = io_b[52 : 0];
  assign adder_adds_1_io_A_1 = io_b[111 : 53];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[53];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[52 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1149 (
  input      [101:0]  io_a,
  input      [101:0]  io_b,
  input               io_c,
  output     [102:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [42:0]   adder_adds_0_io_A_0;
  wire       [42:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [43:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [42:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4139 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[42:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[42:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[43:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[42 : 0];
  assign adder_adds_1_io_A_0 = io_a[101 : 43];
  assign adder_adds_0_io_A_1 = io_b[42 : 0];
  assign adder_adds_1_io_A_1 = io_b[101 : 43];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[43];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[42 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1148 (
  input      [91:0]   io_a,
  input      [91:0]   io_b,
  input               io_c,
  output     [92:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [32:0]   adder_adds_0_io_A_0;
  wire       [32:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [33:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [32:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_4141 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[32:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[32:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[33:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[32 : 0];
  assign adder_adds_1_io_A_0 = io_a[91 : 33];
  assign adder_adds_0_io_A_1 = io_b[32 : 0];
  assign adder_adds_1_io_A_1 = io_b[91 : 33];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[33];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[32 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1147 (
  input      [106:0]  io_a,
  input      [106:0]  io_b,
  input               io_c,
  output     [107:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[106 : 48];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[106 : 48];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1146 (
  input      [136:0]  io_a,
  input      [136:0]  io_b,
  input               io_c,
  output     [137:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [13:0]   adder_adds_0_io_A_0;
  wire       [13:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [14:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [13:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4145 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[13:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[13:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[14:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[13 : 0];
  assign adder_adds_1_io_A_0 = io_a[77 : 14];
  assign adder_adds_2_io_A_0 = io_a[136 : 78];
  assign adder_adds_0_io_A_1 = io_b[13 : 0];
  assign adder_adds_1_io_A_1 = io_b[77 : 14];
  assign adder_adds_2_io_A_1 = io_b[136 : 78];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[14];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[13 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1145 (
  input      [116:0]  io_a,
  input      [116:0]  io_b,
  input               io_c,
  output     [117:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [57:0]   adder_adds_0_io_A_0;
  wire       [57:0]   adder_adds_0_io_A_1;
  wire       [58:0]   adder_adds_1_io_A_0;
  wire       [58:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_0_io_S;
  wire       [59:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg        [57:0]   _zz_io_s_1;
  reg        [58:0]   _zz_io_s_2;

  ADD_5761 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[57:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[57:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[58:0]  )  //o
  );
  ADD_4223 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[57 : 0];
  assign adder_adds_1_io_A_0 = io_a[116 : 58];
  assign adder_adds_0_io_A_1 = io_b[57 : 0];
  assign adder_adds_1_io_A_1 = io_b[116 : 58];
  assign io_s = {_zz_io_s,{_zz_io_s_2,_zz_io_s_1}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[58];
    _zz_io_s <= adder_adds_1_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[57 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[58 : 0];
  end


endmodule

module BADD_1144 (
  input      [154:0]  io_a,
  input      [154:0]  io_b,
  input               io_c,
  output     [155:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [31:0]   adder_adds_0_io_A_0;
  wire       [31:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [32:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [31:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4150 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[31:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[31:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[32:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[31 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 32];
  assign adder_adds_2_io_A_0 = io_a[154 : 96];
  assign adder_adds_0_io_A_1 = io_b[31 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 32];
  assign adder_adds_2_io_A_1 = io_b[154 : 96];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[32];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[31 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1143 (
  input      [262:0]  io_a,
  input      [262:0]  io_b,
  input               io_c,
  output     [263:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [11:0]   adder_adds_0_io_A_0;
  wire       [11:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [58:0]   adder_adds_4_io_A_0;
  wire       [58:0]   adder_adds_4_io_A_1;
  wire       [12:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [59:0]   adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [11:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [58:0]   _zz_io_s_5;

  ADD_4153 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[11:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[11:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[12:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[11 : 0];
  assign adder_adds_1_io_A_0 = io_a[75 : 12];
  assign adder_adds_2_io_A_0 = io_a[139 : 76];
  assign adder_adds_3_io_A_0 = io_a[203 : 140];
  assign adder_adds_4_io_A_0 = io_a[262 : 204];
  assign adder_adds_0_io_A_1 = io_b[11 : 0];
  assign adder_adds_1_io_A_1 = io_b[75 : 12];
  assign adder_adds_2_io_A_1 = io_b[139 : 76];
  assign adder_adds_3_io_A_1 = io_b[203 : 140];
  assign adder_adds_4_io_A_1 = io_b[262 : 204];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[12];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_s <= adder_adds_4_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[11 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[58 : 0];
  end


endmodule

module BADD_1142 (
  input      [214:0]  io_a,
  input      [214:0]  io_b,
  input               io_c,
  output     [215:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [27:0]   adder_adds_0_io_A_0;
  wire       [27:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [28:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [27:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_4158 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[27:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[27:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[28:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[27 : 0];
  assign adder_adds_1_io_A_0 = io_a[91 : 28];
  assign adder_adds_2_io_A_0 = io_a[155 : 92];
  assign adder_adds_3_io_A_0 = io_a[214 : 156];
  assign adder_adds_0_io_A_1 = io_b[27 : 0];
  assign adder_adds_1_io_A_1 = io_b[91 : 28];
  assign adder_adds_2_io_A_1 = io_b[155 : 92];
  assign adder_adds_3_io_A_1 = io_b[214 : 156];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[28];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[27 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1141 (
  input      [176:0]  io_a,
  input      [176:0]  io_b,
  input               io_c,
  output     [177:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [53:0]   adder_adds_0_io_A_0;
  wire       [53:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [54:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [53:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_4162 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[53:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[53:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[54:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[53 : 0];
  assign adder_adds_1_io_A_0 = io_a[117 : 54];
  assign adder_adds_2_io_A_0 = io_a[176 : 118];
  assign adder_adds_0_io_A_1 = io_b[53 : 0];
  assign adder_adds_1_io_A_1 = io_b[117 : 54];
  assign adder_adds_2_io_A_1 = io_b[176 : 118];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[54];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[53 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1140 (
  input      [170:0]  io_a,
  input      [170:0]  io_b,
  input               io_c,
  output     [171:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [58:0]   adder_adds_2_io_A_0;
  wire       [58:0]   adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [59:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [58:0]   _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[111 : 48];
  assign adder_adds_2_io_A_0 = io_a[170 : 112];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[111 : 48];
  assign adder_adds_2_io_A_1 = io_b[170 : 112];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= adder_adds_2_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[58 : 0];
  end


endmodule

module BADD_1139 (
  input      [209:0]  io_a,
  input      [209:0]  io_b,
  input               io_c,
  output     [210:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [22:0]   adder_adds_0_io_A_0;
  wire       [22:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [23:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [22:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_4168 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[22:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[22:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[23:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[22 : 0];
  assign adder_adds_1_io_A_0 = io_a[86 : 23];
  assign adder_adds_2_io_A_0 = io_a[150 : 87];
  assign adder_adds_3_io_A_0 = io_a[209 : 151];
  assign adder_adds_0_io_A_1 = io_b[22 : 0];
  assign adder_adds_1_io_A_1 = io_b[86 : 23];
  assign adder_adds_2_io_A_1 = io_b[150 : 87];
  assign adder_adds_3_io_A_1 = io_b[209 : 151];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[23];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[22 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1138 (
  input      [239:0]  io_a,
  input      [239:0]  io_b,
  input               io_c,
  output     [240:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [52:0]   adder_adds_0_io_A_0;
  wire       [52:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [53:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [52:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_4172 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[52:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[52:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[53:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[52 : 0];
  assign adder_adds_1_io_A_0 = io_a[116 : 53];
  assign adder_adds_2_io_A_0 = io_a[180 : 117];
  assign adder_adds_3_io_A_0 = io_a[239 : 181];
  assign adder_adds_0_io_A_1 = io_b[52 : 0];
  assign adder_adds_1_io_A_1 = io_b[116 : 53];
  assign adder_adds_2_io_A_1 = io_b[180 : 117];
  assign adder_adds_3_io_A_1 = io_b[239 : 181];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[53];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[52 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1137 (
  input      [234:0]  io_a,
  input      [234:0]  io_b,
  input               io_c,
  output     [235:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [58:0]   adder_adds_3_io_A_0;
  wire       [58:0]   adder_adds_3_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [59:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[111 : 48];
  assign adder_adds_2_io_A_0 = io_a[175 : 112];
  assign adder_adds_3_io_A_0 = io_a[234 : 176];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[111 : 48];
  assign adder_adds_2_io_A_1 = io_b[175 : 112];
  assign adder_adds_3_io_A_1 = io_b[234 : 176];
  assign io_s = {_zz_io_s,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_s <= adder_adds_3_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[58 : 0];
  end


endmodule

module BADD_1136 (
  input      [253:0]  io_a,
  input      [253:0]  io_b,
  input               io_c,
  output     [254:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [2:0]    adder_adds_0_io_A_0;
  wire       [2:0]    adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [58:0]   adder_adds_4_io_A_0;
  wire       [58:0]   adder_adds_4_io_A_1;
  wire       [3:0]    adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [59:0]   adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [2:0]    _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [58:0]   _zz_io_s_5;

  ADD_11592 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[2:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[2:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[3:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[2 : 0];
  assign adder_adds_1_io_A_0 = io_a[66 : 3];
  assign adder_adds_2_io_A_0 = io_a[130 : 67];
  assign adder_adds_3_io_A_0 = io_a[194 : 131];
  assign adder_adds_4_io_A_0 = io_a[253 : 195];
  assign adder_adds_0_io_A_1 = io_b[2 : 0];
  assign adder_adds_1_io_A_1 = io_b[66 : 3];
  assign adder_adds_2_io_A_1 = io_b[130 : 67];
  assign adder_adds_3_io_A_1 = io_b[194 : 131];
  assign adder_adds_4_io_A_1 = io_b[253 : 195];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[3];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_s <= adder_adds_4_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[2 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[58 : 0];
  end


endmodule

module BADD_1135 (
  input      [315:0]  io_a,
  input      [315:0]  io_b,
  input               io_c,
  output     [316:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [0:0]    adder_adds_0_io_A_0;
  wire       [0:0]    adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [58:0]   adder_adds_5_io_A_0;
  wire       [58:0]   adder_adds_5_io_A_1;
  wire       [1:0]    adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [59:0]   adder_adds_5_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [0:0]    _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [58:0]   _zz_io_s_6;

  ADD_11601 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0   ), //i
    .io_A_1 (adder_adds_0_io_A_1   ), //i
    .io_CIN (io_c                  ), //i
    .io_S   (adder_adds_0_io_S[1:0])  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[0 : 0];
  assign adder_adds_1_io_A_0 = io_a[64 : 1];
  assign adder_adds_2_io_A_0 = io_a[128 : 65];
  assign adder_adds_3_io_A_0 = io_a[192 : 129];
  assign adder_adds_4_io_A_0 = io_a[256 : 193];
  assign adder_adds_5_io_A_0 = io_a[315 : 257];
  assign adder_adds_0_io_A_1 = io_b[0 : 0];
  assign adder_adds_1_io_A_1 = io_b[64 : 1];
  assign adder_adds_2_io_A_1 = io_b[128 : 65];
  assign adder_adds_3_io_A_1 = io_b[192 : 129];
  assign adder_adds_4_io_A_1 = io_b[256 : 193];
  assign adder_adds_5_io_A_1 = io_b[315 : 257];
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[1];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= adder_adds_5_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[0 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[58 : 0];
  end


endmodule

module BADD_1134 (
  input      [280:0]  io_a,
  input      [280:0]  io_b,
  input               io_c,
  output     [281:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [29:0]   adder_adds_0_io_A_0;
  wire       [29:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [58:0]   adder_adds_4_io_A_0;
  wire       [58:0]   adder_adds_4_io_A_1;
  wire       [30:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [59:0]   adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [29:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [58:0]   _zz_io_s_5;

  ADD_4191 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[29:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[29:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[30:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[29 : 0];
  assign adder_adds_1_io_A_0 = io_a[93 : 30];
  assign adder_adds_2_io_A_0 = io_a[157 : 94];
  assign adder_adds_3_io_A_0 = io_a[221 : 158];
  assign adder_adds_4_io_A_0 = io_a[280 : 222];
  assign adder_adds_0_io_A_1 = io_b[29 : 0];
  assign adder_adds_1_io_A_1 = io_b[93 : 30];
  assign adder_adds_2_io_A_1 = io_b[157 : 94];
  assign adder_adds_3_io_A_1 = io_b[221 : 158];
  assign adder_adds_4_io_A_1 = io_b[280 : 222];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[30];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_s <= adder_adds_4_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[29 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[58 : 0];
  end


endmodule

module BADD_1133 (
  input      [276:0]  io_a,
  input      [276:0]  io_b,
  input               io_c,
  output     [277:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [25:0]   adder_adds_0_io_A_0;
  wire       [25:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [58:0]   adder_adds_4_io_A_0;
  wire       [58:0]   adder_adds_4_io_A_1;
  wire       [26:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [59:0]   adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [25:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [58:0]   _zz_io_s_5;

  ADD_4196 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[25:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[25:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[26:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[25 : 0];
  assign adder_adds_1_io_A_0 = io_a[89 : 26];
  assign adder_adds_2_io_A_0 = io_a[153 : 90];
  assign adder_adds_3_io_A_0 = io_a[217 : 154];
  assign adder_adds_4_io_A_0 = io_a[276 : 218];
  assign adder_adds_0_io_A_1 = io_b[25 : 0];
  assign adder_adds_1_io_A_1 = io_b[89 : 26];
  assign adder_adds_2_io_A_1 = io_b[153 : 90];
  assign adder_adds_3_io_A_1 = io_b[217 : 154];
  assign adder_adds_4_io_A_1 = io_b[276 : 218];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[26];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_s <= adder_adds_4_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[25 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[58 : 0];
  end


endmodule

module BADD_1132 (
  input      [286:0]  io_a,
  input      [286:0]  io_b,
  input               io_c,
  output     [287:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [35:0]   adder_adds_0_io_A_0;
  wire       [35:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [58:0]   adder_adds_4_io_A_0;
  wire       [58:0]   adder_adds_4_io_A_1;
  wire       [36:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [59:0]   adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [35:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [58:0]   _zz_io_s_5;

  ADD_4201 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[35:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[35:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[36:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[35 : 0];
  assign adder_adds_1_io_A_0 = io_a[99 : 36];
  assign adder_adds_2_io_A_0 = io_a[163 : 100];
  assign adder_adds_3_io_A_0 = io_a[227 : 164];
  assign adder_adds_4_io_A_0 = io_a[286 : 228];
  assign adder_adds_0_io_A_1 = io_b[35 : 0];
  assign adder_adds_1_io_A_1 = io_b[99 : 36];
  assign adder_adds_2_io_A_1 = io_b[163 : 100];
  assign adder_adds_3_io_A_1 = io_b[227 : 164];
  assign adder_adds_4_io_A_1 = io_b[286 : 228];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[36];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_s <= adder_adds_4_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[35 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[58 : 0];
  end


endmodule

module BADD_1131 (
  input      [327:0]  io_a,
  input      [327:0]  io_b,
  input               io_c,
  output     [328:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [12:0]   adder_adds_0_io_A_0;
  wire       [12:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [58:0]   adder_adds_5_io_A_0;
  wire       [58:0]   adder_adds_5_io_A_1;
  wire       [13:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [59:0]   adder_adds_5_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [12:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [58:0]   _zz_io_s_6;

  ADD_4237 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[12:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[12:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[13:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[12 : 0];
  assign adder_adds_1_io_A_0 = io_a[76 : 13];
  assign adder_adds_2_io_A_0 = io_a[140 : 77];
  assign adder_adds_3_io_A_0 = io_a[204 : 141];
  assign adder_adds_4_io_A_0 = io_a[268 : 205];
  assign adder_adds_5_io_A_0 = io_a[327 : 269];
  assign adder_adds_0_io_A_1 = io_b[12 : 0];
  assign adder_adds_1_io_A_1 = io_b[76 : 13];
  assign adder_adds_2_io_A_1 = io_b[140 : 77];
  assign adder_adds_3_io_A_1 = io_b[204 : 141];
  assign adder_adds_4_io_A_1 = io_b[268 : 205];
  assign adder_adds_5_io_A_1 = io_b[327 : 269];
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[13];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= adder_adds_5_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[12 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[58 : 0];
  end


endmodule

module BADD_1130 (
  input      [322:0]  io_a,
  input      [322:0]  io_b,
  input               io_c,
  output     [323:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [7:0]    adder_adds_0_io_A_0;
  wire       [7:0]    adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [58:0]   adder_adds_5_io_A_0;
  wire       [58:0]   adder_adds_5_io_A_1;
  wire       [8:0]    adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [59:0]   adder_adds_5_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [7:0]    _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [58:0]   _zz_io_s_6;

  ADD_4212 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[7:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[7:0]), //i
    .io_CIN (io_c                    ), //i
    .io_S   (adder_adds_0_io_S[8:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[7 : 0];
  assign adder_adds_1_io_A_0 = io_a[71 : 8];
  assign adder_adds_2_io_A_0 = io_a[135 : 72];
  assign adder_adds_3_io_A_0 = io_a[199 : 136];
  assign adder_adds_4_io_A_0 = io_a[263 : 200];
  assign adder_adds_5_io_A_0 = io_a[322 : 264];
  assign adder_adds_0_io_A_1 = io_b[7 : 0];
  assign adder_adds_1_io_A_1 = io_b[71 : 8];
  assign adder_adds_2_io_A_1 = io_b[135 : 72];
  assign adder_adds_3_io_A_1 = io_b[199 : 136];
  assign adder_adds_4_io_A_1 = io_b[263 : 200];
  assign adder_adds_5_io_A_1 = io_b[322 : 264];
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[8];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= adder_adds_5_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[7 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[58 : 0];
  end


endmodule

module BADD_1129 (
  input      [332:0]  io_a,
  input      [332:0]  io_b,
  input               io_c,
  output     [333:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [17:0]   adder_adds_0_io_A_0;
  wire       [17:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [58:0]   adder_adds_5_io_A_0;
  wire       [58:0]   adder_adds_5_io_A_1;
  wire       [18:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [59:0]   adder_adds_5_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [17:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [58:0]   _zz_io_s_6;

  ADD_4218 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[17:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[17:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[18:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_4223 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[58:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[58:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[59:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[17 : 0];
  assign adder_adds_1_io_A_0 = io_a[81 : 18];
  assign adder_adds_2_io_A_0 = io_a[145 : 82];
  assign adder_adds_3_io_A_0 = io_a[209 : 146];
  assign adder_adds_4_io_A_0 = io_a[273 : 210];
  assign adder_adds_5_io_A_0 = io_a[332 : 274];
  assign adder_adds_0_io_A_1 = io_b[17 : 0];
  assign adder_adds_1_io_A_1 = io_b[81 : 18];
  assign adder_adds_2_io_A_1 = io_b[145 : 82];
  assign adder_adds_3_io_A_1 = io_b[209 : 146];
  assign adder_adds_4_io_A_1 = io_b[273 : 210];
  assign adder_adds_5_io_A_1 = io_b[332 : 274];
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[18];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= adder_adds_5_io_S[59];
    _zz_io_s_1 <= adder_adds_0_io_S[17 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[58 : 0];
  end


endmodule

module BADD_1128 (
  input      [189:0]  io_a,
  input      [189:0]  io_b,
  input               io_c,
  output     [190:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [61:0]   adder_adds_2_io_A_0;
  wire       [61:0]   adder_adds_2_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [62:0]   adder_adds_2_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [61:0]   _zz_io_A_0_1;
  reg        [61:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_1;
  reg        [61:0]   _zz_io_A_1_1;
  reg        [61:0]   _zz_io_A_1_2;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [61:0]   _zz_io_s_3;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_4226 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[61:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[61:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[62:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_0_io_A_1 = (~ io_b[63 : 0]);
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[189 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_1 <= (~ io_b[127 : 64]);
    _zz_io_A_1_1 <= (~ io_b[189 : 128]);
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_s <= (! adder_adds_2_io_S[62]);
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[61 : 0];
  end


endmodule

module BADD_1127 (
  input      [272:0]  io_a,
  input      [272:0]  io_b,
  input               io_c,
  output     [273:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [16:0]   adder_adds_4_io_A_0;
  wire       [16:0]   adder_adds_4_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [17:0]   adder_adds_4_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [16:0]   _zz_io_A_0_6;
  reg        [16:0]   _zz_io_A_0_7;
  reg        [16:0]   _zz_io_A_0_8;
  reg        [16:0]   _zz_io_A_0_9;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [16:0]   _zz_io_A_1_6;
  reg        [16:0]   _zz_io_A_1_7;
  reg        [16:0]   _zz_io_A_1_8;
  reg        [16:0]   _zz_io_A_1_9;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [16:0]   _zz_io_s_5;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_4231 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[16:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[16:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[17:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_0_io_A_1 = io_b[63 : 0];
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[272 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_1 <= io_b[127 : 64];
    _zz_io_A_1_1 <= io_b[191 : 128];
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= io_b[255 : 192];
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= io_b[272 : 256];
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_s <= adder_adds_4_io_S[17];
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[16 : 0];
  end


endmodule

module BADD_1126 (
  input      [332:0]  io_a,
  input      [332:0]  io_b,
  input               io_c,
  output     [333:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [12:0]   adder_adds_5_io_A_0;
  wire       [12:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [13:0]   adder_adds_5_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [63:0]   _zz_io_A_0_6;
  reg        [63:0]   _zz_io_A_0_7;
  reg        [63:0]   _zz_io_A_0_8;
  reg        [63:0]   _zz_io_A_0_9;
  reg        [12:0]   _zz_io_A_0_10;
  reg        [12:0]   _zz_io_A_0_11;
  reg        [12:0]   _zz_io_A_0_12;
  reg        [12:0]   _zz_io_A_0_13;
  reg        [12:0]   _zz_io_A_0_14;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [63:0]   _zz_io_A_1_6;
  reg        [63:0]   _zz_io_A_1_7;
  reg        [63:0]   _zz_io_A_1_8;
  reg        [63:0]   _zz_io_A_1_9;
  reg        [12:0]   _zz_io_A_1_10;
  reg        [12:0]   _zz_io_A_1_11;
  reg        [12:0]   _zz_io_A_1_12;
  reg        [12:0]   _zz_io_A_1_13;
  reg        [12:0]   _zz_io_A_1_14;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [12:0]   _zz_io_s_6;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_4237 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[12:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[12:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[13:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_5_io_A_0 = _zz_io_A_0_14;
  assign adder_adds_0_io_A_1 = io_b[63 : 0];
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign adder_adds_5_io_A_1 = _zz_io_A_1_14;
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[319 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_0_10 <= io_a[332 : 320];
    _zz_io_A_0_11 <= _zz_io_A_0_10;
    _zz_io_A_0_12 <= _zz_io_A_0_11;
    _zz_io_A_0_13 <= _zz_io_A_0_12;
    _zz_io_A_0_14 <= _zz_io_A_0_13;
    _zz_io_A_1 <= io_b[127 : 64];
    _zz_io_A_1_1 <= io_b[191 : 128];
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= io_b[255 : 192];
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= io_b[319 : 256];
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_A_1_10 <= io_b[332 : 320];
    _zz_io_A_1_11 <= _zz_io_A_1_10;
    _zz_io_A_1_12 <= _zz_io_A_1_11;
    _zz_io_A_1_13 <= _zz_io_A_1_12;
    _zz_io_A_1_14 <= _zz_io_A_1_13;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= adder_adds_5_io_S[13];
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[12 : 0];
  end


endmodule

module BADD_1125 (
  input      [322:0]  io_a,
  input      [322:0]  io_b,
  input               io_c,
  output     [323:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [2:0]    adder_adds_5_io_A_0;
  wire       [2:0]    adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [3:0]    adder_adds_5_io_S;
  reg        [63:0]   _zz_io_A_0;
  reg        [63:0]   _zz_io_A_0_1;
  reg        [63:0]   _zz_io_A_0_2;
  reg        [63:0]   _zz_io_A_0_3;
  reg        [63:0]   _zz_io_A_0_4;
  reg        [63:0]   _zz_io_A_0_5;
  reg        [63:0]   _zz_io_A_0_6;
  reg        [63:0]   _zz_io_A_0_7;
  reg        [63:0]   _zz_io_A_0_8;
  reg        [63:0]   _zz_io_A_0_9;
  reg        [2:0]    _zz_io_A_0_10;
  reg        [2:0]    _zz_io_A_0_11;
  reg        [2:0]    _zz_io_A_0_12;
  reg        [2:0]    _zz_io_A_0_13;
  reg        [2:0]    _zz_io_A_0_14;
  reg        [63:0]   _zz_io_A_1;
  reg        [63:0]   _zz_io_A_1_1;
  reg        [63:0]   _zz_io_A_1_2;
  reg        [63:0]   _zz_io_A_1_3;
  reg        [63:0]   _zz_io_A_1_4;
  reg        [63:0]   _zz_io_A_1_5;
  reg        [63:0]   _zz_io_A_1_6;
  reg        [63:0]   _zz_io_A_1_7;
  reg        [63:0]   _zz_io_A_1_8;
  reg        [63:0]   _zz_io_A_1_9;
  reg        [2:0]    _zz_io_A_1_10;
  reg        [2:0]    _zz_io_A_1_11;
  reg        [2:0]    _zz_io_A_1_12;
  reg        [2:0]    _zz_io_A_1_13;
  reg        [2:0]    _zz_io_A_1_14;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [2:0]    _zz_io_s_6;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_11592 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[2:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[2:0]), //i
    .io_CIN (_zz_io_CIN_4            ), //i
    .io_S   (adder_adds_5_io_S[3:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = _zz_io_A_0;
  assign adder_adds_2_io_A_0 = _zz_io_A_0_2;
  assign adder_adds_3_io_A_0 = _zz_io_A_0_5;
  assign adder_adds_4_io_A_0 = _zz_io_A_0_9;
  assign adder_adds_5_io_A_0 = _zz_io_A_0_14;
  assign adder_adds_0_io_A_1 = io_b[63 : 0];
  assign adder_adds_1_io_A_1 = _zz_io_A_1;
  assign adder_adds_2_io_A_1 = _zz_io_A_1_2;
  assign adder_adds_3_io_A_1 = _zz_io_A_1_5;
  assign adder_adds_4_io_A_1 = _zz_io_A_1_9;
  assign adder_adds_5_io_A_1 = _zz_io_A_1_14;
  assign io_s = {_zz_io_s,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}};
  always @(posedge clk) begin
    _zz_io_A_0 <= io_a[127 : 64];
    _zz_io_A_0_1 <= io_a[191 : 128];
    _zz_io_A_0_2 <= _zz_io_A_0_1;
    _zz_io_A_0_3 <= io_a[255 : 192];
    _zz_io_A_0_4 <= _zz_io_A_0_3;
    _zz_io_A_0_5 <= _zz_io_A_0_4;
    _zz_io_A_0_6 <= io_a[319 : 256];
    _zz_io_A_0_7 <= _zz_io_A_0_6;
    _zz_io_A_0_8 <= _zz_io_A_0_7;
    _zz_io_A_0_9 <= _zz_io_A_0_8;
    _zz_io_A_0_10 <= io_a[322 : 320];
    _zz_io_A_0_11 <= _zz_io_A_0_10;
    _zz_io_A_0_12 <= _zz_io_A_0_11;
    _zz_io_A_0_13 <= _zz_io_A_0_12;
    _zz_io_A_0_14 <= _zz_io_A_0_13;
    _zz_io_A_1 <= io_b[127 : 64];
    _zz_io_A_1_1 <= io_b[191 : 128];
    _zz_io_A_1_2 <= _zz_io_A_1_1;
    _zz_io_A_1_3 <= io_b[255 : 192];
    _zz_io_A_1_4 <= _zz_io_A_1_3;
    _zz_io_A_1_5 <= _zz_io_A_1_4;
    _zz_io_A_1_6 <= io_b[319 : 256];
    _zz_io_A_1_7 <= _zz_io_A_1_6;
    _zz_io_A_1_8 <= _zz_io_A_1_7;
    _zz_io_A_1_9 <= _zz_io_A_1_8;
    _zz_io_A_1_10 <= io_b[322 : 320];
    _zz_io_A_1_11 <= _zz_io_A_1_10;
    _zz_io_A_1_12 <= _zz_io_A_1_11;
    _zz_io_A_1_13 <= _zz_io_A_1_12;
    _zz_io_A_1_14 <= _zz_io_A_1_13;
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= adder_adds_5_io_S[3];
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[2 : 0];
  end


endmodule

//KaratsubaCore_34 replaced by KaratsubaCore_35

module KaratsubaCore_35 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_a_2,
  input      [47:0]   io_a_3,
  input      [47:0]   io_a_4,
  input      [47:0]   io_a_5,
  input      [47:0]   io_a_6,
  input      [47:0]   io_a_7,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  input      [47:0]   io_b_2,
  input      [47:0]   io_b_3,
  input      [47:0]   io_b_4,
  input      [47:0]   io_b_5,
  input      [47:0]   io_b_6,
  input      [47:0]   io_b_7,
  output reg [767:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [384:0]  karatsuba_add2_io_a;
  wire       [575:0]  karatsuba_noExtend_add3_io_a;
  reg        [575:0]  karatsuba_noExtend_add3_io_b;
  wire       [383:0]  karatsuba_lsbMul_io_p;
  wire       [385:0]  karatsuba_midMul_io_p;
  wire       [383:0]  karatsuba_msbMul_io_p;
  wire       [48:0]   karatsuba_midAdd_0_0_io_S;
  wire       [48:0]   karatsuba_midAdd_0_1_io_S;
  wire       [48:0]   karatsuba_midAdd_0_2_io_S;
  wire       [48:0]   karatsuba_midAdd_0_3_io_S;
  wire       [48:0]   karatsuba_midAdd_1_0_io_S;
  wire       [48:0]   karatsuba_midAdd_1_1_io_S;
  wire       [48:0]   karatsuba_midAdd_1_2_io_S;
  wire       [48:0]   karatsuba_midAdd_1_3_io_S;
  wire       [384:0]  karatsuba_add1_io_s;
  wire       [385:0]  karatsuba_add2_io_s;
  wire       [576:0]  karatsuba_noExtend_add3_io_s;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_a_1;
  reg        [48:0]   _zz_io_a_2;
  reg        [48:0]   _zz_io_a_3;
  reg        [48:0]   _zz_io_b_0;
  reg        [48:0]   _zz_io_b_1;
  reg        [48:0]   _zz_io_b_2;
  reg        [48:0]   _zz_io_b_3;
  reg        [384:0]  core_karatsuba_add1_io_s_delay_1;
  reg        [384:0]  _zz_io_a;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_1;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_2;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_3;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_4;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_5;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_6;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_7;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_8;
  reg        [191:0]  _zz_io_p;

  KaratsubaCore_141 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]                ), //i
    .io_a_1 (io_a_1[47:0]                ), //i
    .io_a_2 (io_a_2[47:0]                ), //i
    .io_a_3 (io_a_3[47:0]                ), //i
    .io_b_0 (io_b_0[47:0]                ), //i
    .io_b_1 (io_b_1[47:0]                ), //i
    .io_b_2 (io_b_2[47:0]                ), //i
    .io_b_3 (io_b_3[47:0]                ), //i
    .io_p   (karatsuba_lsbMul_io_p[383:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_142 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]            ), //i
    .io_a_1 (_zz_io_a_1[48:0]            ), //i
    .io_a_2 (_zz_io_a_2[48:0]            ), //i
    .io_a_3 (_zz_io_a_3[48:0]            ), //i
    .io_b_0 (_zz_io_b_0[48:0]            ), //i
    .io_b_1 (_zz_io_b_1[48:0]            ), //i
    .io_b_2 (_zz_io_b_2[48:0]            ), //i
    .io_b_3 (_zz_io_b_3[48:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[385:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_143 karatsuba_msbMul (
    .io_a_0 (io_a_4[47:0]                ), //i
    .io_a_1 (io_a_5[47:0]                ), //i
    .io_a_2 (io_a_6[47:0]                ), //i
    .io_a_3 (io_a_7[47:0]                ), //i
    .io_b_0 (io_b_4[47:0]                ), //i
    .io_b_1 (io_b_5[47:0]                ), //i
    .io_b_2 (io_b_6[47:0]                ), //i
    .io_b_3 (io_b_7[47:0]                ), //i
    .io_p   (karatsuba_msbMul_io_p[383:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  ADD_11602 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[47:0]                   ), //i
    .io_A_1 (io_a_4[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_0_1 (
    .io_A_0 (io_a_1[47:0]                   ), //i
    .io_A_1 (io_a_5[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_1_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_0_2 (
    .io_A_0 (io_a_2[47:0]                   ), //i
    .io_A_1 (io_a_6[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_2_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_0_3 (
    .io_A_0 (io_a_3[47:0]                   ), //i
    .io_A_1 (io_a_7[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_3_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[47:0]                   ), //i
    .io_A_1 (io_b_4[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_1 (
    .io_A_0 (io_b_1[47:0]                   ), //i
    .io_A_1 (io_b_5[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_1_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_2 (
    .io_A_0 (io_b_2[47:0]                   ), //i
    .io_A_1 (io_b_6[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_2_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_3 (
    .io_A_0 (io_b_3[47:0]                   ), //i
    .io_A_1 (io_b_7[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_3_io_S[48:0])  //o
  );
  BADD_1310 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[383:0]), //i
    .io_b   (karatsuba_msbMul_io_p[383:0]), //i
    .io_c   (1'b0                        ), //i
    .io_s   (karatsuba_add1_io_s[384:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_1311 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[384:0]             ), //i
    .io_b   (core_karatsuba_add1_io_s_delay_1[384:0]), //i
    .io_c   (1'b1                                   ), //i
    .io_s   (karatsuba_add2_io_s[385:0]             ), //o
    .clk    (clk                                    ), //i
    .resetn (resetn                                 )  //i
  );
  BADD_1312 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[575:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[575:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[576:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[384:0];
  assign karatsuba_noExtend_add3_io_a = {191'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[191 : 0] = (karatsuba_lsbMul_io_p >>> 192);
    karatsuba_noExtend_add3_io_b[575 : 192] = core_karatsuba_msbMul_io_p_delay_8;
  end

  always @(*) begin
    io_p[191 : 0] = _zz_io_p;
    io_p[767 : 192] = karatsuba_noExtend_add3_io_s[575:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_a_1 <= karatsuba_midAdd_0_1_io_S;
    _zz_io_a_2 <= karatsuba_midAdd_0_2_io_S;
    _zz_io_a_3 <= karatsuba_midAdd_0_3_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b_1 <= karatsuba_midAdd_1_1_io_S;
    _zz_io_b_2 <= karatsuba_midAdd_1_2_io_S;
    _zz_io_b_3 <= karatsuba_midAdd_1_3_io_S;
    core_karatsuba_add1_io_s_delay_1 <= karatsuba_add1_io_s;
    _zz_io_a <= karatsuba_add2_io_s[384:0];
    core_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    core_karatsuba_msbMul_io_p_delay_2 <= core_karatsuba_msbMul_io_p_delay_1;
    core_karatsuba_msbMul_io_p_delay_3 <= core_karatsuba_msbMul_io_p_delay_2;
    core_karatsuba_msbMul_io_p_delay_4 <= core_karatsuba_msbMul_io_p_delay_3;
    core_karatsuba_msbMul_io_p_delay_5 <= core_karatsuba_msbMul_io_p_delay_4;
    core_karatsuba_msbMul_io_p_delay_6 <= core_karatsuba_msbMul_io_p_delay_5;
    core_karatsuba_msbMul_io_p_delay_7 <= core_karatsuba_msbMul_io_p_delay_6;
    core_karatsuba_msbMul_io_p_delay_8 <= core_karatsuba_msbMul_io_p_delay_7;
    _zz_io_p <= karatsuba_lsbMul_io_p[191 : 0];
  end


endmodule

//ADD_227 replaced by ADD_5761

//ADD_226 replaced by ADD_5756

//ADD_225 replaced by ADD_5756

//ADD_224 replaced by ADD_5756

//ADD_223 replaced by ADD_5756

//ADD_222 replaced by ADD_5756

//ADD_233 replaced by ADD_5761

//ADD_232 replaced by ADD_5756

//ADD_231 replaced by ADD_5756

//ADD_230 replaced by ADD_5756

//ADD_229 replaced by ADD_5756

//ADD_228 replaced by ADD_5756

//ADD_239 replaced by ADD_5761

//ADD_238 replaced by ADD_5756

//ADD_237 replaced by ADD_5756

//ADD_236 replaced by ADD_5756

//ADD_235 replaced by ADD_5756

//ADD_234 replaced by ADD_5756

//ADD_245 replaced by ADD_5761

//ADD_244 replaced by ADD_5756

//ADD_243 replaced by ADD_5756

//ADD_242 replaced by ADD_5756

//ADD_241 replaced by ADD_5756

//ADD_240 replaced by ADD_5756

//ADD_251 replaced by ADD_5761

//ADD_250 replaced by ADD_5756

//ADD_249 replaced by ADD_5756

//ADD_248 replaced by ADD_5756

//ADD_247 replaced by ADD_5756

//ADD_246 replaced by ADD_5756

//ADD_257 replaced by ADD_5761

//ADD_256 replaced by ADD_5756

//ADD_255 replaced by ADD_5756

//ADD_254 replaced by ADD_5756

//ADD_253 replaced by ADD_5756

//ADD_252 replaced by ADD_5756

//ADD_263 replaced by ADD_5761

//ADD_262 replaced by ADD_5756

//ADD_261 replaced by ADD_5756

//ADD_260 replaced by ADD_5756

//ADD_259 replaced by ADD_5756

//ADD_258 replaced by ADD_5756

//ADD_269 replaced by ADD_5761

//ADD_268 replaced by ADD_5756

//ADD_267 replaced by ADD_5756

//ADD_266 replaced by ADD_5756

//ADD_265 replaced by ADD_5756

//ADD_264 replaced by ADD_5756

//BADD_1187 replaced by BADD_1306

//ADD_275 replaced by ADD_5761

//ADD_274 replaced by ADD_5756

//ADD_273 replaced by ADD_5756

//ADD_272 replaced by ADD_5756

//ADD_271 replaced by ADD_5756

//ADD_270 replaced by ADD_5756

//ADD_281 replaced by ADD_4223

//ADD_280 replaced by ADD_5756

//ADD_279 replaced by ADD_5756

//ADD_278 replaced by ADD_5756

//ADD_277 replaced by ADD_5756

//ADD_276 replaced by ADD_5756

//ADD_283 replaced by ADD_4223

//ADD_282 replaced by ADD_4226

//ADD_284 replaced by ADD_4055

//ADD_285 replaced by ADD_4057

//ADD_287 replaced by ADD_4223

//ADD_286 replaced by ADD_4057

//ADD_288 replaced by ADD_4223

//ADD_289 replaced by ADD_4060

//ADD_291 replaced by ADD_4223

//ADD_290 replaced by ADD_11560

//ADD_293 replaced by ADD_4223

//ADD_292 replaced by ADD_4196

//ADD_295 replaced by ADD_4223

//ADD_294 replaced by ADD_4132

//ADD_297 replaced by ADD_4223

//ADD_296 replaced by ADD_4067

//ADD_301 replaced by ADD_4223

//ADD_300 replaced by ADD_5756

//ADD_299 replaced by ADD_5756

//ADD_298 replaced by ADD_11592

//ADD_304 replaced by ADD_4223

//ADD_303 replaced by ADD_5756

//ADD_302 replaced by ADD_4168

//ADD_307 replaced by ADD_4223

//ADD_306 replaced by ADD_5756

//ADD_305 replaced by ADD_4076

//ADD_310 replaced by ADD_4223

//ADD_309 replaced by ADD_5756

//ADD_308 replaced by ADD_11592

//ADD_313 replaced by ADD_4223

//ADD_312 replaced by ADD_5756

//ADD_311 replaced by ADD_4106

//ADD_316 replaced by ADD_4223

//ADD_315 replaced by ADD_5756

//ADD_314 replaced by ADD_4085

//ADD_319 replaced by ADD_4223

//ADD_318 replaced by ADD_5756

//ADD_317 replaced by ADD_4158

//ADD_322 replaced by ADD_4223

//ADD_321 replaced by ADD_5756

//ADD_320 replaced by ADD_4091

//ADD_326 replaced by ADD_4223

//ADD_325 replaced by ADD_5756

//ADD_324 replaced by ADD_5756

//ADD_323 replaced by ADD_4094

//ADD_330 replaced by ADD_4223

//ADD_329 replaced by ADD_5756

//ADD_328 replaced by ADD_5756

//ADD_327 replaced by ADD_4145

//ADD_334 replaced by ADD_4223

//ADD_333 replaced by ADD_5756

//ADD_332 replaced by ADD_5756

//ADD_331 replaced by ADD_4212

//ADD_338 replaced by ADD_4223

//ADD_337 replaced by ADD_5756

//ADD_336 replaced by ADD_5756

//ADD_335 replaced by ADD_4106

//ADD_343 replaced by ADD_4223

//ADD_342 replaced by ADD_5756

//ADD_341 replaced by ADD_5756

//ADD_340 replaced by ADD_5756

//ADD_339 replaced by ADD_4212

//ADD_347 replaced by ADD_4223

//ADD_346 replaced by ADD_5756

//ADD_345 replaced by ADD_5756

//ADD_344 replaced by ADD_4115

//ADD_352 replaced by ADD_4223

//ADD_351 replaced by ADD_5756

//ADD_350 replaced by ADD_5756

//ADD_349 replaced by ADD_5756

//ADD_348 replaced by ADD_4231

//ADD_353 replaced by ADD_11560

//ADD_356 replaced by ADD_4223

//ADD_355 replaced by ADD_5756

//ADD_354 replaced by ADD_4125

//ADD_358 replaced by ADD_4223

//ADD_357 replaced by ADD_4131

//ADD_359 replaced by ADD_4150

//ADD_360 replaced by ADD_4131

//ADD_361 replaced by ADD_4132

//ADD_362 replaced by ADD_4196

//ADD_363 replaced by ADD_4134

//ADD_364 replaced by ADD_4139

//ADD_365 replaced by ADD_4136

//ADD_367 replaced by ADD_4223

//ADD_366 replaced by ADD_4172

//ADD_369 replaced by ADD_4223

//ADD_368 replaced by ADD_4139

//ADD_371 replaced by ADD_4223

//ADD_370 replaced by ADD_4141

//ADD_373 replaced by ADD_4223

//ADD_372 replaced by ADD_11602

//ADD_376 replaced by ADD_4223

//ADD_375 replaced by ADD_5756

//ADD_374 replaced by ADD_4145

//ADD_378 replaced by ADD_4223

//ADD_377 replaced by ADD_5761

//ADD_381 replaced by ADD_4223

//ADD_380 replaced by ADD_5756

//ADD_379 replaced by ADD_4150

//ADD_386 replaced by ADD_4223

//ADD_385 replaced by ADD_5756

//ADD_384 replaced by ADD_5756

//ADD_383 replaced by ADD_5756

//ADD_382 replaced by ADD_4153

//ADD_390 replaced by ADD_4223

//ADD_389 replaced by ADD_5756

//ADD_388 replaced by ADD_5756

//ADD_387 replaced by ADD_4158

//ADD_393 replaced by ADD_4223

//ADD_392 replaced by ADD_5756

//ADD_391 replaced by ADD_4162

//ADD_396 replaced by ADD_4223

//ADD_395 replaced by ADD_5756

//ADD_394 replaced by ADD_11602

//ADD_400 replaced by ADD_4223

//ADD_399 replaced by ADD_5756

//ADD_398 replaced by ADD_5756

//ADD_397 replaced by ADD_4168

//ADD_404 replaced by ADD_4223

//ADD_403 replaced by ADD_5756

//ADD_402 replaced by ADD_5756

//ADD_401 replaced by ADD_4172

//ADD_408 replaced by ADD_4223

//ADD_407 replaced by ADD_5756

//ADD_406 replaced by ADD_5756

//ADD_405 replaced by ADD_11602

//ADD_413 replaced by ADD_4223

//ADD_412 replaced by ADD_5756

//ADD_411 replaced by ADD_5756

//ADD_410 replaced by ADD_5756

//ADD_409 replaced by ADD_11592

//ADD_419 replaced by ADD_4223

//ADD_418 replaced by ADD_5756

//ADD_417 replaced by ADD_5756

//ADD_416 replaced by ADD_5756

//ADD_415 replaced by ADD_5756

//ADD_414 replaced by ADD_11601

//ADD_424 replaced by ADD_4223

//ADD_423 replaced by ADD_5756

//ADD_422 replaced by ADD_5756

//ADD_421 replaced by ADD_5756

//ADD_420 replaced by ADD_4191

//ADD_429 replaced by ADD_4223

//ADD_428 replaced by ADD_5756

//ADD_427 replaced by ADD_5756

//ADD_426 replaced by ADD_5756

//ADD_425 replaced by ADD_4196

//ADD_434 replaced by ADD_4223

//ADD_433 replaced by ADD_5756

//ADD_432 replaced by ADD_5756

//ADD_431 replaced by ADD_5756

//ADD_430 replaced by ADD_4201

//ADD_440 replaced by ADD_4223

//ADD_439 replaced by ADD_5756

//ADD_438 replaced by ADD_5756

//ADD_437 replaced by ADD_5756

//ADD_436 replaced by ADD_5756

//ADD_435 replaced by ADD_4237

//ADD_446 replaced by ADD_4223

//ADD_445 replaced by ADD_5756

//ADD_444 replaced by ADD_5756

//ADD_443 replaced by ADD_5756

//ADD_442 replaced by ADD_5756

//ADD_441 replaced by ADD_4212

//ADD_452 replaced by ADD_4223

//ADD_451 replaced by ADD_5756

//ADD_450 replaced by ADD_5756

//ADD_449 replaced by ADD_5756

//ADD_448 replaced by ADD_5756

//ADD_447 replaced by ADD_4218

//ADD_455 replaced by ADD_4226

//ADD_454 replaced by ADD_5756

//ADD_453 replaced by ADD_5756

//ADD_460 replaced by ADD_4231

//ADD_459 replaced by ADD_5756

//ADD_458 replaced by ADD_5756

//ADD_457 replaced by ADD_5756

//ADD_456 replaced by ADD_5756

//ADD_466 replaced by ADD_4237

//ADD_465 replaced by ADD_5756

//ADD_464 replaced by ADD_5756

//ADD_463 replaced by ADD_5756

//ADD_462 replaced by ADD_5756

//ADD_461 replaced by ADD_5756

//ADD_472 replaced by ADD_11592

//ADD_471 replaced by ADD_5756

//ADD_470 replaced by ADD_5756

//ADD_469 replaced by ADD_5756

//ADD_468 replaced by ADD_5756

//ADD_467 replaced by ADD_5756

//BADD_1190 replaced by BADD_1312

//BADD_1189 replaced by BADD_1311

//BADD_1188 replaced by BADD_1310

//ADD_480 replaced by ADD_11602

//ADD_479 replaced by ADD_11602

//ADD_478 replaced by ADD_11602

//ADD_477 replaced by ADD_11602

//ADD_476 replaced by ADD_11602

//ADD_475 replaced by ADD_11602

//ADD_474 replaced by ADD_11602

//ADD_473 replaced by ADD_11602

//KaratsubaCore_38 replaced by KaratsubaCore_143

//KaratsubaCore_37 replaced by KaratsubaCore_142

//KaratsubaCore_36 replaced by KaratsubaCore_141

//BADD_1193 replaced by BADD_1312

//BADD_1192 replaced by BADD_1311

//BADD_1191 replaced by BADD_1310

//ADD_488 replaced by ADD_11602

//ADD_487 replaced by ADD_11602

//ADD_486 replaced by ADD_11602

//ADD_485 replaced by ADD_11602

//ADD_484 replaced by ADD_11602

//ADD_483 replaced by ADD_11602

//ADD_482 replaced by ADD_11602

//ADD_481 replaced by ADD_11602

//KaratsubaCore_41 replaced by KaratsubaCore_143

//KaratsubaCore_40 replaced by KaratsubaCore_142

//KaratsubaCore_39 replaced by KaratsubaCore_141

//BADD_1194 replaced by BADD_1306

//ADD_494 replaced by ADD_5761

//ADD_493 replaced by ADD_5756

//ADD_492 replaced by ADD_5756

//ADD_491 replaced by ADD_5756

//ADD_490 replaced by ADD_5756

//ADD_489 replaced by ADD_5756

//ADD_500 replaced by ADD_4223

//ADD_499 replaced by ADD_5756

//ADD_498 replaced by ADD_5756

//ADD_497 replaced by ADD_5756

//ADD_496 replaced by ADD_5756

//ADD_495 replaced by ADD_5756

//ADD_502 replaced by ADD_4223

//ADD_501 replaced by ADD_4226

//ADD_503 replaced by ADD_4055

//ADD_504 replaced by ADD_4057

//ADD_506 replaced by ADD_4223

//ADD_505 replaced by ADD_4057

//ADD_507 replaced by ADD_4223

//ADD_508 replaced by ADD_4060

//ADD_510 replaced by ADD_4223

//ADD_509 replaced by ADD_11560

//ADD_512 replaced by ADD_4223

//ADD_511 replaced by ADD_4196

//ADD_514 replaced by ADD_4223

//ADD_513 replaced by ADD_4132

//ADD_516 replaced by ADD_4223

//ADD_515 replaced by ADD_4067

//ADD_520 replaced by ADD_4223

//ADD_519 replaced by ADD_5756

//ADD_518 replaced by ADD_5756

//ADD_517 replaced by ADD_11592

//ADD_523 replaced by ADD_4223

//ADD_522 replaced by ADD_5756

//ADD_521 replaced by ADD_4168

//ADD_526 replaced by ADD_4223

//ADD_525 replaced by ADD_5756

//ADD_524 replaced by ADD_4076

//ADD_529 replaced by ADD_4223

//ADD_528 replaced by ADD_5756

//ADD_527 replaced by ADD_11592

//ADD_532 replaced by ADD_4223

//ADD_531 replaced by ADD_5756

//ADD_530 replaced by ADD_4106

//ADD_535 replaced by ADD_4223

//ADD_534 replaced by ADD_5756

//ADD_533 replaced by ADD_4085

//ADD_538 replaced by ADD_4223

//ADD_537 replaced by ADD_5756

//ADD_536 replaced by ADD_4158

//ADD_541 replaced by ADD_4223

//ADD_540 replaced by ADD_5756

//ADD_539 replaced by ADD_4091

//ADD_545 replaced by ADD_4223

//ADD_544 replaced by ADD_5756

//ADD_543 replaced by ADD_5756

//ADD_542 replaced by ADD_4094

//ADD_549 replaced by ADD_4223

//ADD_548 replaced by ADD_5756

//ADD_547 replaced by ADD_5756

//ADD_546 replaced by ADD_4145

//ADD_553 replaced by ADD_4223

//ADD_552 replaced by ADD_5756

//ADD_551 replaced by ADD_5756

//ADD_550 replaced by ADD_4212

//ADD_557 replaced by ADD_4223

//ADD_556 replaced by ADD_5756

//ADD_555 replaced by ADD_5756

//ADD_554 replaced by ADD_4106

//ADD_562 replaced by ADD_4223

//ADD_561 replaced by ADD_5756

//ADD_560 replaced by ADD_5756

//ADD_559 replaced by ADD_5756

//ADD_558 replaced by ADD_4212

//ADD_566 replaced by ADD_4223

//ADD_565 replaced by ADD_5756

//ADD_564 replaced by ADD_5756

//ADD_563 replaced by ADD_4115

//ADD_571 replaced by ADD_4223

//ADD_570 replaced by ADD_5756

//ADD_569 replaced by ADD_5756

//ADD_568 replaced by ADD_5756

//ADD_567 replaced by ADD_4231

//ADD_572 replaced by ADD_11560

//ADD_575 replaced by ADD_4223

//ADD_574 replaced by ADD_5756

//ADD_573 replaced by ADD_4125

//ADD_577 replaced by ADD_4223

//ADD_576 replaced by ADD_4131

//ADD_578 replaced by ADD_4150

//ADD_579 replaced by ADD_4131

//ADD_580 replaced by ADD_4132

//ADD_581 replaced by ADD_4196

//ADD_582 replaced by ADD_4134

//ADD_583 replaced by ADD_4139

//ADD_584 replaced by ADD_4136

//ADD_586 replaced by ADD_4223

//ADD_585 replaced by ADD_4172

//ADD_588 replaced by ADD_4223

//ADD_587 replaced by ADD_4139

//ADD_590 replaced by ADD_4223

//ADD_589 replaced by ADD_4141

//ADD_592 replaced by ADD_4223

//ADD_591 replaced by ADD_11602

//ADD_595 replaced by ADD_4223

//ADD_594 replaced by ADD_5756

//ADD_593 replaced by ADD_4145

//ADD_597 replaced by ADD_4223

//ADD_596 replaced by ADD_5761

//ADD_600 replaced by ADD_4223

//ADD_599 replaced by ADD_5756

//ADD_598 replaced by ADD_4150

//ADD_605 replaced by ADD_4223

//ADD_604 replaced by ADD_5756

//ADD_603 replaced by ADD_5756

//ADD_602 replaced by ADD_5756

//ADD_601 replaced by ADD_4153

//ADD_609 replaced by ADD_4223

//ADD_608 replaced by ADD_5756

//ADD_607 replaced by ADD_5756

//ADD_606 replaced by ADD_4158

//ADD_612 replaced by ADD_4223

//ADD_611 replaced by ADD_5756

//ADD_610 replaced by ADD_4162

//ADD_615 replaced by ADD_4223

//ADD_614 replaced by ADD_5756

//ADD_613 replaced by ADD_11602

//ADD_619 replaced by ADD_4223

//ADD_618 replaced by ADD_5756

//ADD_617 replaced by ADD_5756

//ADD_616 replaced by ADD_4168

//ADD_623 replaced by ADD_4223

//ADD_622 replaced by ADD_5756

//ADD_621 replaced by ADD_5756

//ADD_620 replaced by ADD_4172

//ADD_627 replaced by ADD_4223

//ADD_626 replaced by ADD_5756

//ADD_625 replaced by ADD_5756

//ADD_624 replaced by ADD_11602

//ADD_632 replaced by ADD_4223

//ADD_631 replaced by ADD_5756

//ADD_630 replaced by ADD_5756

//ADD_629 replaced by ADD_5756

//ADD_628 replaced by ADD_11592

//ADD_638 replaced by ADD_4223

//ADD_637 replaced by ADD_5756

//ADD_636 replaced by ADD_5756

//ADD_635 replaced by ADD_5756

//ADD_634 replaced by ADD_5756

//ADD_633 replaced by ADD_11601

//ADD_643 replaced by ADD_4223

//ADD_642 replaced by ADD_5756

//ADD_641 replaced by ADD_5756

//ADD_640 replaced by ADD_5756

//ADD_639 replaced by ADD_4191

//ADD_648 replaced by ADD_4223

//ADD_647 replaced by ADD_5756

//ADD_646 replaced by ADD_5756

//ADD_645 replaced by ADD_5756

//ADD_644 replaced by ADD_4196

//ADD_653 replaced by ADD_4223

//ADD_652 replaced by ADD_5756

//ADD_651 replaced by ADD_5756

//ADD_650 replaced by ADD_5756

//ADD_649 replaced by ADD_4201

//ADD_659 replaced by ADD_4223

//ADD_658 replaced by ADD_5756

//ADD_657 replaced by ADD_5756

//ADD_656 replaced by ADD_5756

//ADD_655 replaced by ADD_5756

//ADD_654 replaced by ADD_4237

//ADD_665 replaced by ADD_4223

//ADD_664 replaced by ADD_5756

//ADD_663 replaced by ADD_5756

//ADD_662 replaced by ADD_5756

//ADD_661 replaced by ADD_5756

//ADD_660 replaced by ADD_4212

//ADD_671 replaced by ADD_4223

//ADD_670 replaced by ADD_5756

//ADD_669 replaced by ADD_5756

//ADD_668 replaced by ADD_5756

//ADD_667 replaced by ADD_5756

//ADD_666 replaced by ADD_4218

//ADD_674 replaced by ADD_4226

//ADD_673 replaced by ADD_5756

//ADD_672 replaced by ADD_5756

//ADD_679 replaced by ADD_4231

//ADD_678 replaced by ADD_5756

//ADD_677 replaced by ADD_5756

//ADD_676 replaced by ADD_5756

//ADD_675 replaced by ADD_5756

//ADD_685 replaced by ADD_4237

//ADD_684 replaced by ADD_5756

//ADD_683 replaced by ADD_5756

//ADD_682 replaced by ADD_5756

//ADD_681 replaced by ADD_5756

//ADD_680 replaced by ADD_5756

//ADD_691 replaced by ADD_11592

//ADD_690 replaced by ADD_5756

//ADD_689 replaced by ADD_5756

//ADD_688 replaced by ADD_5756

//ADD_687 replaced by ADD_5756

//ADD_686 replaced by ADD_5756

//BADD_1197 replaced by BADD_1312

//BADD_1196 replaced by BADD_1311

//BADD_1195 replaced by BADD_1310

//ADD_699 replaced by ADD_11602

//ADD_698 replaced by ADD_11602

//ADD_697 replaced by ADD_11602

//ADD_696 replaced by ADD_11602

//ADD_695 replaced by ADD_11602

//ADD_694 replaced by ADD_11602

//ADD_693 replaced by ADD_11602

//ADD_692 replaced by ADD_11602

//KaratsubaCore_44 replaced by KaratsubaCore_143

//KaratsubaCore_43 replaced by KaratsubaCore_142

//KaratsubaCore_42 replaced by KaratsubaCore_141

//BADD_1200 replaced by BADD_1312

//BADD_1199 replaced by BADD_1311

//BADD_1198 replaced by BADD_1310

//ADD_707 replaced by ADD_11602

//ADD_706 replaced by ADD_11602

//ADD_705 replaced by ADD_11602

//ADD_704 replaced by ADD_11602

//ADD_703 replaced by ADD_11602

//ADD_702 replaced by ADD_11602

//ADD_701 replaced by ADD_11602

//ADD_700 replaced by ADD_11602

//KaratsubaCore_47 replaced by KaratsubaCore_143

//KaratsubaCore_46 replaced by KaratsubaCore_142

//KaratsubaCore_45 replaced by KaratsubaCore_141

//BADD_1201 replaced by BADD_1306

//ADD_713 replaced by ADD_5761

//ADD_712 replaced by ADD_5756

//ADD_711 replaced by ADD_5756

//ADD_710 replaced by ADD_5756

//ADD_709 replaced by ADD_5756

//ADD_708 replaced by ADD_5756

//ADD_719 replaced by ADD_4223

//ADD_718 replaced by ADD_5756

//ADD_717 replaced by ADD_5756

//ADD_716 replaced by ADD_5756

//ADD_715 replaced by ADD_5756

//ADD_714 replaced by ADD_5756

//ADD_721 replaced by ADD_4223

//ADD_720 replaced by ADD_4226

//ADD_722 replaced by ADD_4055

//ADD_723 replaced by ADD_4057

//ADD_725 replaced by ADD_4223

//ADD_724 replaced by ADD_4057

//ADD_726 replaced by ADD_4223

//ADD_727 replaced by ADD_4060

//ADD_729 replaced by ADD_4223

//ADD_728 replaced by ADD_11560

//ADD_731 replaced by ADD_4223

//ADD_730 replaced by ADD_4196

//ADD_733 replaced by ADD_4223

//ADD_732 replaced by ADD_4132

//ADD_735 replaced by ADD_4223

//ADD_734 replaced by ADD_4067

//ADD_739 replaced by ADD_4223

//ADD_738 replaced by ADD_5756

//ADD_737 replaced by ADD_5756

//ADD_736 replaced by ADD_11592

//ADD_742 replaced by ADD_4223

//ADD_741 replaced by ADD_5756

//ADD_740 replaced by ADD_4168

//ADD_745 replaced by ADD_4223

//ADD_744 replaced by ADD_5756

//ADD_743 replaced by ADD_4076

//ADD_748 replaced by ADD_4223

//ADD_747 replaced by ADD_5756

//ADD_746 replaced by ADD_11592

//ADD_751 replaced by ADD_4223

//ADD_750 replaced by ADD_5756

//ADD_749 replaced by ADD_4106

//ADD_754 replaced by ADD_4223

//ADD_753 replaced by ADD_5756

//ADD_752 replaced by ADD_4085

//ADD_757 replaced by ADD_4223

//ADD_756 replaced by ADD_5756

//ADD_755 replaced by ADD_4158

//ADD_760 replaced by ADD_4223

//ADD_759 replaced by ADD_5756

//ADD_758 replaced by ADD_4091

//ADD_764 replaced by ADD_4223

//ADD_763 replaced by ADD_5756

//ADD_762 replaced by ADD_5756

//ADD_761 replaced by ADD_4094

//ADD_768 replaced by ADD_4223

//ADD_767 replaced by ADD_5756

//ADD_766 replaced by ADD_5756

//ADD_765 replaced by ADD_4145

//ADD_772 replaced by ADD_4223

//ADD_771 replaced by ADD_5756

//ADD_770 replaced by ADD_5756

//ADD_769 replaced by ADD_4212

//ADD_776 replaced by ADD_4223

//ADD_775 replaced by ADD_5756

//ADD_774 replaced by ADD_5756

//ADD_773 replaced by ADD_4106

//ADD_781 replaced by ADD_4223

//ADD_780 replaced by ADD_5756

//ADD_779 replaced by ADD_5756

//ADD_778 replaced by ADD_5756

//ADD_777 replaced by ADD_4212

//ADD_785 replaced by ADD_4223

//ADD_784 replaced by ADD_5756

//ADD_783 replaced by ADD_5756

//ADD_782 replaced by ADD_4115

//ADD_790 replaced by ADD_4223

//ADD_789 replaced by ADD_5756

//ADD_788 replaced by ADD_5756

//ADD_787 replaced by ADD_5756

//ADD_786 replaced by ADD_4231

//ADD_791 replaced by ADD_11560

//ADD_794 replaced by ADD_4223

//ADD_793 replaced by ADD_5756

//ADD_792 replaced by ADD_4125

//ADD_796 replaced by ADD_4223

//ADD_795 replaced by ADD_4131

//ADD_797 replaced by ADD_4150

//ADD_798 replaced by ADD_4131

//ADD_799 replaced by ADD_4132

//ADD_800 replaced by ADD_4196

//ADD_801 replaced by ADD_4134

//ADD_802 replaced by ADD_4139

//ADD_803 replaced by ADD_4136

//ADD_805 replaced by ADD_4223

//ADD_804 replaced by ADD_4172

//ADD_807 replaced by ADD_4223

//ADD_806 replaced by ADD_4139

//ADD_809 replaced by ADD_4223

//ADD_808 replaced by ADD_4141

//ADD_811 replaced by ADD_4223

//ADD_810 replaced by ADD_11602

//ADD_814 replaced by ADD_4223

//ADD_813 replaced by ADD_5756

//ADD_812 replaced by ADD_4145

//ADD_816 replaced by ADD_4223

//ADD_815 replaced by ADD_5761

//ADD_819 replaced by ADD_4223

//ADD_818 replaced by ADD_5756

//ADD_817 replaced by ADD_4150

//ADD_824 replaced by ADD_4223

//ADD_823 replaced by ADD_5756

//ADD_822 replaced by ADD_5756

//ADD_821 replaced by ADD_5756

//ADD_820 replaced by ADD_4153

//ADD_828 replaced by ADD_4223

//ADD_827 replaced by ADD_5756

//ADD_826 replaced by ADD_5756

//ADD_825 replaced by ADD_4158

//ADD_831 replaced by ADD_4223

//ADD_830 replaced by ADD_5756

//ADD_829 replaced by ADD_4162

//ADD_834 replaced by ADD_4223

//ADD_833 replaced by ADD_5756

//ADD_832 replaced by ADD_11602

//ADD_838 replaced by ADD_4223

//ADD_837 replaced by ADD_5756

//ADD_836 replaced by ADD_5756

//ADD_835 replaced by ADD_4168

//ADD_842 replaced by ADD_4223

//ADD_841 replaced by ADD_5756

//ADD_840 replaced by ADD_5756

//ADD_839 replaced by ADD_4172

//ADD_846 replaced by ADD_4223

//ADD_845 replaced by ADD_5756

//ADD_844 replaced by ADD_5756

//ADD_843 replaced by ADD_11602

//ADD_851 replaced by ADD_4223

//ADD_850 replaced by ADD_5756

//ADD_849 replaced by ADD_5756

//ADD_848 replaced by ADD_5756

//ADD_847 replaced by ADD_11592

//ADD_857 replaced by ADD_4223

//ADD_856 replaced by ADD_5756

//ADD_855 replaced by ADD_5756

//ADD_854 replaced by ADD_5756

//ADD_853 replaced by ADD_5756

//ADD_852 replaced by ADD_11601

//ADD_862 replaced by ADD_4223

//ADD_861 replaced by ADD_5756

//ADD_860 replaced by ADD_5756

//ADD_859 replaced by ADD_5756

//ADD_858 replaced by ADD_4191

//ADD_867 replaced by ADD_4223

//ADD_866 replaced by ADD_5756

//ADD_865 replaced by ADD_5756

//ADD_864 replaced by ADD_5756

//ADD_863 replaced by ADD_4196

//ADD_872 replaced by ADD_4223

//ADD_871 replaced by ADD_5756

//ADD_870 replaced by ADD_5756

//ADD_869 replaced by ADD_5756

//ADD_868 replaced by ADD_4201

//ADD_878 replaced by ADD_4223

//ADD_877 replaced by ADD_5756

//ADD_876 replaced by ADD_5756

//ADD_875 replaced by ADD_5756

//ADD_874 replaced by ADD_5756

//ADD_873 replaced by ADD_4237

//ADD_884 replaced by ADD_4223

//ADD_883 replaced by ADD_5756

//ADD_882 replaced by ADD_5756

//ADD_881 replaced by ADD_5756

//ADD_880 replaced by ADD_5756

//ADD_879 replaced by ADD_4212

//ADD_890 replaced by ADD_4223

//ADD_889 replaced by ADD_5756

//ADD_888 replaced by ADD_5756

//ADD_887 replaced by ADD_5756

//ADD_886 replaced by ADD_5756

//ADD_885 replaced by ADD_4218

//ADD_893 replaced by ADD_4226

//ADD_892 replaced by ADD_5756

//ADD_891 replaced by ADD_5756

//ADD_898 replaced by ADD_4231

//ADD_897 replaced by ADD_5756

//ADD_896 replaced by ADD_5756

//ADD_895 replaced by ADD_5756

//ADD_894 replaced by ADD_5756

//ADD_904 replaced by ADD_4237

//ADD_903 replaced by ADD_5756

//ADD_902 replaced by ADD_5756

//ADD_901 replaced by ADD_5756

//ADD_900 replaced by ADD_5756

//ADD_899 replaced by ADD_5756

//ADD_910 replaced by ADD_11592

//ADD_909 replaced by ADD_5756

//ADD_908 replaced by ADD_5756

//ADD_907 replaced by ADD_5756

//ADD_906 replaced by ADD_5756

//ADD_905 replaced by ADD_5756

//BADD_1204 replaced by BADD_1312

//BADD_1203 replaced by BADD_1311

//BADD_1202 replaced by BADD_1310

//ADD_918 replaced by ADD_11602

//ADD_917 replaced by ADD_11602

//ADD_916 replaced by ADD_11602

//ADD_915 replaced by ADD_11602

//ADD_914 replaced by ADD_11602

//ADD_913 replaced by ADD_11602

//ADD_912 replaced by ADD_11602

//ADD_911 replaced by ADD_11602

//KaratsubaCore_50 replaced by KaratsubaCore_143

//KaratsubaCore_49 replaced by KaratsubaCore_142

//KaratsubaCore_48 replaced by KaratsubaCore_141

//BADD_1207 replaced by BADD_1312

//BADD_1206 replaced by BADD_1311

//BADD_1205 replaced by BADD_1310

//ADD_926 replaced by ADD_11602

//ADD_925 replaced by ADD_11602

//ADD_924 replaced by ADD_11602

//ADD_923 replaced by ADD_11602

//ADD_922 replaced by ADD_11602

//ADD_921 replaced by ADD_11602

//ADD_920 replaced by ADD_11602

//ADD_919 replaced by ADD_11602

//KaratsubaCore_53 replaced by KaratsubaCore_143

//KaratsubaCore_52 replaced by KaratsubaCore_142

//KaratsubaCore_51 replaced by KaratsubaCore_141

//BADD_1208 replaced by BADD_1306

//ADD_932 replaced by ADD_5761

//ADD_931 replaced by ADD_5756

//ADD_930 replaced by ADD_5756

//ADD_929 replaced by ADD_5756

//ADD_928 replaced by ADD_5756

//ADD_927 replaced by ADD_5756

//ADD_938 replaced by ADD_4223

//ADD_937 replaced by ADD_5756

//ADD_936 replaced by ADD_5756

//ADD_935 replaced by ADD_5756

//ADD_934 replaced by ADD_5756

//ADD_933 replaced by ADD_5756

//ADD_940 replaced by ADD_4223

//ADD_939 replaced by ADD_4226

//ADD_941 replaced by ADD_4055

//ADD_942 replaced by ADD_4057

//ADD_944 replaced by ADD_4223

//ADD_943 replaced by ADD_4057

//ADD_945 replaced by ADD_4223

//ADD_946 replaced by ADD_4060

//ADD_948 replaced by ADD_4223

//ADD_947 replaced by ADD_11560

//ADD_950 replaced by ADD_4223

//ADD_949 replaced by ADD_4196

//ADD_952 replaced by ADD_4223

//ADD_951 replaced by ADD_4132

//ADD_954 replaced by ADD_4223

//ADD_953 replaced by ADD_4067

//ADD_958 replaced by ADD_4223

//ADD_957 replaced by ADD_5756

//ADD_956 replaced by ADD_5756

//ADD_955 replaced by ADD_11592

//ADD_961 replaced by ADD_4223

//ADD_960 replaced by ADD_5756

//ADD_959 replaced by ADD_4168

//ADD_964 replaced by ADD_4223

//ADD_963 replaced by ADD_5756

//ADD_962 replaced by ADD_4076

//ADD_967 replaced by ADD_4223

//ADD_966 replaced by ADD_5756

//ADD_965 replaced by ADD_11592

//ADD_970 replaced by ADD_4223

//ADD_969 replaced by ADD_5756

//ADD_968 replaced by ADD_4106

//ADD_973 replaced by ADD_4223

//ADD_972 replaced by ADD_5756

//ADD_971 replaced by ADD_4085

//ADD_976 replaced by ADD_4223

//ADD_975 replaced by ADD_5756

//ADD_974 replaced by ADD_4158

//ADD_979 replaced by ADD_4223

//ADD_978 replaced by ADD_5756

//ADD_977 replaced by ADD_4091

//ADD_983 replaced by ADD_4223

//ADD_982 replaced by ADD_5756

//ADD_981 replaced by ADD_5756

//ADD_980 replaced by ADD_4094

//ADD_987 replaced by ADD_4223

//ADD_986 replaced by ADD_5756

//ADD_985 replaced by ADD_5756

//ADD_984 replaced by ADD_4145

//ADD_991 replaced by ADD_4223

//ADD_990 replaced by ADD_5756

//ADD_989 replaced by ADD_5756

//ADD_988 replaced by ADD_4212

//ADD_995 replaced by ADD_4223

//ADD_994 replaced by ADD_5756

//ADD_993 replaced by ADD_5756

//ADD_992 replaced by ADD_4106

//ADD_1000 replaced by ADD_4223

//ADD_999 replaced by ADD_5756

//ADD_998 replaced by ADD_5756

//ADD_997 replaced by ADD_5756

//ADD_996 replaced by ADD_4212

//ADD_1004 replaced by ADD_4223

//ADD_1003 replaced by ADD_5756

//ADD_1002 replaced by ADD_5756

//ADD_1001 replaced by ADD_4115

//ADD_1009 replaced by ADD_4223

//ADD_1008 replaced by ADD_5756

//ADD_1007 replaced by ADD_5756

//ADD_1006 replaced by ADD_5756

//ADD_1005 replaced by ADD_4231

//ADD_1010 replaced by ADD_11560

//ADD_1013 replaced by ADD_4223

//ADD_1012 replaced by ADD_5756

//ADD_1011 replaced by ADD_4125

//ADD_1015 replaced by ADD_4223

//ADD_1014 replaced by ADD_4131

//ADD_1016 replaced by ADD_4150

//ADD_1017 replaced by ADD_4131

//ADD_1018 replaced by ADD_4132

//ADD_1019 replaced by ADD_4196

//ADD_1020 replaced by ADD_4134

//ADD_1021 replaced by ADD_4139

//ADD_1022 replaced by ADD_4136

//ADD_1024 replaced by ADD_4223

//ADD_1023 replaced by ADD_4172

//ADD_1026 replaced by ADD_4223

//ADD_1025 replaced by ADD_4139

//ADD_1028 replaced by ADD_4223

//ADD_1027 replaced by ADD_4141

//ADD_1030 replaced by ADD_4223

//ADD_1029 replaced by ADD_11602

//ADD_1033 replaced by ADD_4223

//ADD_1032 replaced by ADD_5756

//ADD_1031 replaced by ADD_4145

//ADD_1035 replaced by ADD_4223

//ADD_1034 replaced by ADD_5761

//ADD_1038 replaced by ADD_4223

//ADD_1037 replaced by ADD_5756

//ADD_1036 replaced by ADD_4150

//ADD_1043 replaced by ADD_4223

//ADD_1042 replaced by ADD_5756

//ADD_1041 replaced by ADD_5756

//ADD_1040 replaced by ADD_5756

//ADD_1039 replaced by ADD_4153

//ADD_1047 replaced by ADD_4223

//ADD_1046 replaced by ADD_5756

//ADD_1045 replaced by ADD_5756

//ADD_1044 replaced by ADD_4158

//ADD_1050 replaced by ADD_4223

//ADD_1049 replaced by ADD_5756

//ADD_1048 replaced by ADD_4162

//ADD_1053 replaced by ADD_4223

//ADD_1052 replaced by ADD_5756

//ADD_1051 replaced by ADD_11602

//ADD_1057 replaced by ADD_4223

//ADD_1056 replaced by ADD_5756

//ADD_1055 replaced by ADD_5756

//ADD_1054 replaced by ADD_4168

//ADD_1061 replaced by ADD_4223

//ADD_1060 replaced by ADD_5756

//ADD_1059 replaced by ADD_5756

//ADD_1058 replaced by ADD_4172

//ADD_1065 replaced by ADD_4223

//ADD_1064 replaced by ADD_5756

//ADD_1063 replaced by ADD_5756

//ADD_1062 replaced by ADD_11602

//ADD_1070 replaced by ADD_4223

//ADD_1069 replaced by ADD_5756

//ADD_1068 replaced by ADD_5756

//ADD_1067 replaced by ADD_5756

//ADD_1066 replaced by ADD_11592

//ADD_1076 replaced by ADD_4223

//ADD_1075 replaced by ADD_5756

//ADD_1074 replaced by ADD_5756

//ADD_1073 replaced by ADD_5756

//ADD_1072 replaced by ADD_5756

//ADD_1071 replaced by ADD_11601

//ADD_1081 replaced by ADD_4223

//ADD_1080 replaced by ADD_5756

//ADD_1079 replaced by ADD_5756

//ADD_1078 replaced by ADD_5756

//ADD_1077 replaced by ADD_4191

//ADD_1086 replaced by ADD_4223

//ADD_1085 replaced by ADD_5756

//ADD_1084 replaced by ADD_5756

//ADD_1083 replaced by ADD_5756

//ADD_1082 replaced by ADD_4196

//ADD_1091 replaced by ADD_4223

//ADD_1090 replaced by ADD_5756

//ADD_1089 replaced by ADD_5756

//ADD_1088 replaced by ADD_5756

//ADD_1087 replaced by ADD_4201

//ADD_1097 replaced by ADD_4223

//ADD_1096 replaced by ADD_5756

//ADD_1095 replaced by ADD_5756

//ADD_1094 replaced by ADD_5756

//ADD_1093 replaced by ADD_5756

//ADD_1092 replaced by ADD_4237

//ADD_1103 replaced by ADD_4223

//ADD_1102 replaced by ADD_5756

//ADD_1101 replaced by ADD_5756

//ADD_1100 replaced by ADD_5756

//ADD_1099 replaced by ADD_5756

//ADD_1098 replaced by ADD_4212

//ADD_1109 replaced by ADD_4223

//ADD_1108 replaced by ADD_5756

//ADD_1107 replaced by ADD_5756

//ADD_1106 replaced by ADD_5756

//ADD_1105 replaced by ADD_5756

//ADD_1104 replaced by ADD_4218

//ADD_1112 replaced by ADD_4226

//ADD_1111 replaced by ADD_5756

//ADD_1110 replaced by ADD_5756

//ADD_1117 replaced by ADD_4231

//ADD_1116 replaced by ADD_5756

//ADD_1115 replaced by ADD_5756

//ADD_1114 replaced by ADD_5756

//ADD_1113 replaced by ADD_5756

//ADD_1123 replaced by ADD_4237

//ADD_1122 replaced by ADD_5756

//ADD_1121 replaced by ADD_5756

//ADD_1120 replaced by ADD_5756

//ADD_1119 replaced by ADD_5756

//ADD_1118 replaced by ADD_5756

//ADD_1129 replaced by ADD_11592

//ADD_1128 replaced by ADD_5756

//ADD_1127 replaced by ADD_5756

//ADD_1126 replaced by ADD_5756

//ADD_1125 replaced by ADD_5756

//ADD_1124 replaced by ADD_5756

//BADD_1211 replaced by BADD_1312

//BADD_1210 replaced by BADD_1311

//BADD_1209 replaced by BADD_1310

//ADD_1137 replaced by ADD_11602

//ADD_1136 replaced by ADD_11602

//ADD_1135 replaced by ADD_11602

//ADD_1134 replaced by ADD_11602

//ADD_1133 replaced by ADD_11602

//ADD_1132 replaced by ADD_11602

//ADD_1131 replaced by ADD_11602

//ADD_1130 replaced by ADD_11602

//KaratsubaCore_56 replaced by KaratsubaCore_143

//KaratsubaCore_55 replaced by KaratsubaCore_142

//KaratsubaCore_54 replaced by KaratsubaCore_141

//BADD_1214 replaced by BADD_1312

//BADD_1213 replaced by BADD_1311

//BADD_1212 replaced by BADD_1310

//ADD_1145 replaced by ADD_11602

//ADD_1144 replaced by ADD_11602

//ADD_1143 replaced by ADD_11602

//ADD_1142 replaced by ADD_11602

//ADD_1141 replaced by ADD_11602

//ADD_1140 replaced by ADD_11602

//ADD_1139 replaced by ADD_11602

//ADD_1138 replaced by ADD_11602

//KaratsubaCore_59 replaced by KaratsubaCore_143

//KaratsubaCore_58 replaced by KaratsubaCore_142

//KaratsubaCore_57 replaced by KaratsubaCore_141

//BADD_1215 replaced by BADD_1306

//ADD_1151 replaced by ADD_5761

//ADD_1150 replaced by ADD_5756

//ADD_1149 replaced by ADD_5756

//ADD_1148 replaced by ADD_5756

//ADD_1147 replaced by ADD_5756

//ADD_1146 replaced by ADD_5756

//ADD_1157 replaced by ADD_4223

//ADD_1156 replaced by ADD_5756

//ADD_1155 replaced by ADD_5756

//ADD_1154 replaced by ADD_5756

//ADD_1153 replaced by ADD_5756

//ADD_1152 replaced by ADD_5756

//ADD_1159 replaced by ADD_4223

//ADD_1158 replaced by ADD_4226

//ADD_1160 replaced by ADD_4055

//ADD_1161 replaced by ADD_4057

//ADD_1163 replaced by ADD_4223

//ADD_1162 replaced by ADD_4057

//ADD_1164 replaced by ADD_4223

//ADD_1165 replaced by ADD_4060

//ADD_1167 replaced by ADD_4223

//ADD_1166 replaced by ADD_11560

//ADD_1169 replaced by ADD_4223

//ADD_1168 replaced by ADD_4196

//ADD_1171 replaced by ADD_4223

//ADD_1170 replaced by ADD_4132

//ADD_1173 replaced by ADD_4223

//ADD_1172 replaced by ADD_4067

//ADD_1177 replaced by ADD_4223

//ADD_1176 replaced by ADD_5756

//ADD_1175 replaced by ADD_5756

//ADD_1174 replaced by ADD_11592

//ADD_1180 replaced by ADD_4223

//ADD_1179 replaced by ADD_5756

//ADD_1178 replaced by ADD_4168

//ADD_1183 replaced by ADD_4223

//ADD_1182 replaced by ADD_5756

//ADD_1181 replaced by ADD_4076

//ADD_1186 replaced by ADD_4223

//ADD_1185 replaced by ADD_5756

//ADD_1184 replaced by ADD_11592

//ADD_1189 replaced by ADD_4223

//ADD_1188 replaced by ADD_5756

//ADD_1187 replaced by ADD_4106

//ADD_1192 replaced by ADD_4223

//ADD_1191 replaced by ADD_5756

//ADD_1190 replaced by ADD_4085

//ADD_1195 replaced by ADD_4223

//ADD_1194 replaced by ADD_5756

//ADD_1193 replaced by ADD_4158

//ADD_1198 replaced by ADD_4223

//ADD_1197 replaced by ADD_5756

//ADD_1196 replaced by ADD_4091

//ADD_1202 replaced by ADD_4223

//ADD_1201 replaced by ADD_5756

//ADD_1200 replaced by ADD_5756

//ADD_1199 replaced by ADD_4094

//ADD_1206 replaced by ADD_4223

//ADD_1205 replaced by ADD_5756

//ADD_1204 replaced by ADD_5756

//ADD_1203 replaced by ADD_4145

//ADD_1210 replaced by ADD_4223

//ADD_1209 replaced by ADD_5756

//ADD_1208 replaced by ADD_5756

//ADD_1207 replaced by ADD_4212

//ADD_1214 replaced by ADD_4223

//ADD_1213 replaced by ADD_5756

//ADD_1212 replaced by ADD_5756

//ADD_1211 replaced by ADD_4106

//ADD_1219 replaced by ADD_4223

//ADD_1218 replaced by ADD_5756

//ADD_1217 replaced by ADD_5756

//ADD_1216 replaced by ADD_5756

//ADD_1215 replaced by ADD_4212

//ADD_1223 replaced by ADD_4223

//ADD_1222 replaced by ADD_5756

//ADD_1221 replaced by ADD_5756

//ADD_1220 replaced by ADD_4115

//ADD_1228 replaced by ADD_4223

//ADD_1227 replaced by ADD_5756

//ADD_1226 replaced by ADD_5756

//ADD_1225 replaced by ADD_5756

//ADD_1224 replaced by ADD_4231

//ADD_1229 replaced by ADD_11560

//ADD_1232 replaced by ADD_4223

//ADD_1231 replaced by ADD_5756

//ADD_1230 replaced by ADD_4125

//ADD_1234 replaced by ADD_4223

//ADD_1233 replaced by ADD_4131

//ADD_1235 replaced by ADD_4150

//ADD_1236 replaced by ADD_4131

//ADD_1237 replaced by ADD_4132

//ADD_1238 replaced by ADD_4196

//ADD_1239 replaced by ADD_4134

//ADD_1240 replaced by ADD_4139

//ADD_1241 replaced by ADD_4136

//ADD_1243 replaced by ADD_4223

//ADD_1242 replaced by ADD_4172

//ADD_1245 replaced by ADD_4223

//ADD_1244 replaced by ADD_4139

//ADD_1247 replaced by ADD_4223

//ADD_1246 replaced by ADD_4141

//ADD_1249 replaced by ADD_4223

//ADD_1248 replaced by ADD_11602

//ADD_1252 replaced by ADD_4223

//ADD_1251 replaced by ADD_5756

//ADD_1250 replaced by ADD_4145

//ADD_1254 replaced by ADD_4223

//ADD_1253 replaced by ADD_5761

//ADD_1257 replaced by ADD_4223

//ADD_1256 replaced by ADD_5756

//ADD_1255 replaced by ADD_4150

//ADD_1262 replaced by ADD_4223

//ADD_1261 replaced by ADD_5756

//ADD_1260 replaced by ADD_5756

//ADD_1259 replaced by ADD_5756

//ADD_1258 replaced by ADD_4153

//ADD_1266 replaced by ADD_4223

//ADD_1265 replaced by ADD_5756

//ADD_1264 replaced by ADD_5756

//ADD_1263 replaced by ADD_4158

//ADD_1269 replaced by ADD_4223

//ADD_1268 replaced by ADD_5756

//ADD_1267 replaced by ADD_4162

//ADD_1272 replaced by ADD_4223

//ADD_1271 replaced by ADD_5756

//ADD_1270 replaced by ADD_11602

//ADD_1276 replaced by ADD_4223

//ADD_1275 replaced by ADD_5756

//ADD_1274 replaced by ADD_5756

//ADD_1273 replaced by ADD_4168

//ADD_1280 replaced by ADD_4223

//ADD_1279 replaced by ADD_5756

//ADD_1278 replaced by ADD_5756

//ADD_1277 replaced by ADD_4172

//ADD_1284 replaced by ADD_4223

//ADD_1283 replaced by ADD_5756

//ADD_1282 replaced by ADD_5756

//ADD_1281 replaced by ADD_11602

//ADD_1289 replaced by ADD_4223

//ADD_1288 replaced by ADD_5756

//ADD_1287 replaced by ADD_5756

//ADD_1286 replaced by ADD_5756

//ADD_1285 replaced by ADD_11592

//ADD_1295 replaced by ADD_4223

//ADD_1294 replaced by ADD_5756

//ADD_1293 replaced by ADD_5756

//ADD_1292 replaced by ADD_5756

//ADD_1291 replaced by ADD_5756

//ADD_1290 replaced by ADD_11601

//ADD_1300 replaced by ADD_4223

//ADD_1299 replaced by ADD_5756

//ADD_1298 replaced by ADD_5756

//ADD_1297 replaced by ADD_5756

//ADD_1296 replaced by ADD_4191

//ADD_1305 replaced by ADD_4223

//ADD_1304 replaced by ADD_5756

//ADD_1303 replaced by ADD_5756

//ADD_1302 replaced by ADD_5756

//ADD_1301 replaced by ADD_4196

//ADD_1310 replaced by ADD_4223

//ADD_1309 replaced by ADD_5756

//ADD_1308 replaced by ADD_5756

//ADD_1307 replaced by ADD_5756

//ADD_1306 replaced by ADD_4201

//ADD_1316 replaced by ADD_4223

//ADD_1315 replaced by ADD_5756

//ADD_1314 replaced by ADD_5756

//ADD_1313 replaced by ADD_5756

//ADD_1312 replaced by ADD_5756

//ADD_1311 replaced by ADD_4237

//ADD_1322 replaced by ADD_4223

//ADD_1321 replaced by ADD_5756

//ADD_1320 replaced by ADD_5756

//ADD_1319 replaced by ADD_5756

//ADD_1318 replaced by ADD_5756

//ADD_1317 replaced by ADD_4212

//ADD_1328 replaced by ADD_4223

//ADD_1327 replaced by ADD_5756

//ADD_1326 replaced by ADD_5756

//ADD_1325 replaced by ADD_5756

//ADD_1324 replaced by ADD_5756

//ADD_1323 replaced by ADD_4218

//ADD_1331 replaced by ADD_4226

//ADD_1330 replaced by ADD_5756

//ADD_1329 replaced by ADD_5756

//ADD_1336 replaced by ADD_4231

//ADD_1335 replaced by ADD_5756

//ADD_1334 replaced by ADD_5756

//ADD_1333 replaced by ADD_5756

//ADD_1332 replaced by ADD_5756

//ADD_1342 replaced by ADD_4237

//ADD_1341 replaced by ADD_5756

//ADD_1340 replaced by ADD_5756

//ADD_1339 replaced by ADD_5756

//ADD_1338 replaced by ADD_5756

//ADD_1337 replaced by ADD_5756

//ADD_1348 replaced by ADD_11592

//ADD_1347 replaced by ADD_5756

//ADD_1346 replaced by ADD_5756

//ADD_1345 replaced by ADD_5756

//ADD_1344 replaced by ADD_5756

//ADD_1343 replaced by ADD_5756

//BADD_1218 replaced by BADD_1312

//BADD_1217 replaced by BADD_1311

//BADD_1216 replaced by BADD_1310

//ADD_1356 replaced by ADD_11602

//ADD_1355 replaced by ADD_11602

//ADD_1354 replaced by ADD_11602

//ADD_1353 replaced by ADD_11602

//ADD_1352 replaced by ADD_11602

//ADD_1351 replaced by ADD_11602

//ADD_1350 replaced by ADD_11602

//ADD_1349 replaced by ADD_11602

//KaratsubaCore_62 replaced by KaratsubaCore_143

//KaratsubaCore_61 replaced by KaratsubaCore_142

//KaratsubaCore_60 replaced by KaratsubaCore_141

//BADD_1221 replaced by BADD_1312

//BADD_1220 replaced by BADD_1311

//BADD_1219 replaced by BADD_1310

//ADD_1364 replaced by ADD_11602

//ADD_1363 replaced by ADD_11602

//ADD_1362 replaced by ADD_11602

//ADD_1361 replaced by ADD_11602

//ADD_1360 replaced by ADD_11602

//ADD_1359 replaced by ADD_11602

//ADD_1358 replaced by ADD_11602

//ADD_1357 replaced by ADD_11602

//KaratsubaCore_65 replaced by KaratsubaCore_143

//KaratsubaCore_64 replaced by KaratsubaCore_142

//KaratsubaCore_63 replaced by KaratsubaCore_141

//BADD_1222 replaced by BADD_1306

//ADD_1370 replaced by ADD_5761

//ADD_1369 replaced by ADD_5756

//ADD_1368 replaced by ADD_5756

//ADD_1367 replaced by ADD_5756

//ADD_1366 replaced by ADD_5756

//ADD_1365 replaced by ADD_5756

//ADD_1376 replaced by ADD_4223

//ADD_1375 replaced by ADD_5756

//ADD_1374 replaced by ADD_5756

//ADD_1373 replaced by ADD_5756

//ADD_1372 replaced by ADD_5756

//ADD_1371 replaced by ADD_5756

//ADD_1378 replaced by ADD_4223

//ADD_1377 replaced by ADD_4226

//ADD_1379 replaced by ADD_4055

//ADD_1380 replaced by ADD_4057

//ADD_1382 replaced by ADD_4223

//ADD_1381 replaced by ADD_4057

//ADD_1383 replaced by ADD_4223

//ADD_1384 replaced by ADD_4060

//ADD_1386 replaced by ADD_4223

//ADD_1385 replaced by ADD_11560

//ADD_1388 replaced by ADD_4223

//ADD_1387 replaced by ADD_4196

//ADD_1390 replaced by ADD_4223

//ADD_1389 replaced by ADD_4132

//ADD_1392 replaced by ADD_4223

//ADD_1391 replaced by ADD_4067

//ADD_1396 replaced by ADD_4223

//ADD_1395 replaced by ADD_5756

//ADD_1394 replaced by ADD_5756

//ADD_1393 replaced by ADD_11592

//ADD_1399 replaced by ADD_4223

//ADD_1398 replaced by ADD_5756

//ADD_1397 replaced by ADD_4168

//ADD_1402 replaced by ADD_4223

//ADD_1401 replaced by ADD_5756

//ADD_1400 replaced by ADD_4076

//ADD_1405 replaced by ADD_4223

//ADD_1404 replaced by ADD_5756

//ADD_1403 replaced by ADD_11592

//ADD_1408 replaced by ADD_4223

//ADD_1407 replaced by ADD_5756

//ADD_1406 replaced by ADD_4106

//ADD_1411 replaced by ADD_4223

//ADD_1410 replaced by ADD_5756

//ADD_1409 replaced by ADD_4085

//ADD_1414 replaced by ADD_4223

//ADD_1413 replaced by ADD_5756

//ADD_1412 replaced by ADD_4158

//ADD_1417 replaced by ADD_4223

//ADD_1416 replaced by ADD_5756

//ADD_1415 replaced by ADD_4091

//ADD_1421 replaced by ADD_4223

//ADD_1420 replaced by ADD_5756

//ADD_1419 replaced by ADD_5756

//ADD_1418 replaced by ADD_4094

//ADD_1425 replaced by ADD_4223

//ADD_1424 replaced by ADD_5756

//ADD_1423 replaced by ADD_5756

//ADD_1422 replaced by ADD_4145

//ADD_1429 replaced by ADD_4223

//ADD_1428 replaced by ADD_5756

//ADD_1427 replaced by ADD_5756

//ADD_1426 replaced by ADD_4212

//ADD_1433 replaced by ADD_4223

//ADD_1432 replaced by ADD_5756

//ADD_1431 replaced by ADD_5756

//ADD_1430 replaced by ADD_4106

//ADD_1438 replaced by ADD_4223

//ADD_1437 replaced by ADD_5756

//ADD_1436 replaced by ADD_5756

//ADD_1435 replaced by ADD_5756

//ADD_1434 replaced by ADD_4212

//ADD_1442 replaced by ADD_4223

//ADD_1441 replaced by ADD_5756

//ADD_1440 replaced by ADD_5756

//ADD_1439 replaced by ADD_4115

//ADD_1447 replaced by ADD_4223

//ADD_1446 replaced by ADD_5756

//ADD_1445 replaced by ADD_5756

//ADD_1444 replaced by ADD_5756

//ADD_1443 replaced by ADD_4231

//ADD_1448 replaced by ADD_11560

//ADD_1451 replaced by ADD_4223

//ADD_1450 replaced by ADD_5756

//ADD_1449 replaced by ADD_4125

//ADD_1453 replaced by ADD_4223

//ADD_1452 replaced by ADD_4131

//ADD_1454 replaced by ADD_4150

//ADD_1455 replaced by ADD_4131

//ADD_1456 replaced by ADD_4132

//ADD_1457 replaced by ADD_4196

//ADD_1458 replaced by ADD_4134

//ADD_1459 replaced by ADD_4139

//ADD_1460 replaced by ADD_4136

//ADD_1462 replaced by ADD_4223

//ADD_1461 replaced by ADD_4172

//ADD_1464 replaced by ADD_4223

//ADD_1463 replaced by ADD_4139

//ADD_1466 replaced by ADD_4223

//ADD_1465 replaced by ADD_4141

//ADD_1468 replaced by ADD_4223

//ADD_1467 replaced by ADD_11602

//ADD_1471 replaced by ADD_4223

//ADD_1470 replaced by ADD_5756

//ADD_1469 replaced by ADD_4145

//ADD_1473 replaced by ADD_4223

//ADD_1472 replaced by ADD_5761

//ADD_1476 replaced by ADD_4223

//ADD_1475 replaced by ADD_5756

//ADD_1474 replaced by ADD_4150

//ADD_1481 replaced by ADD_4223

//ADD_1480 replaced by ADD_5756

//ADD_1479 replaced by ADD_5756

//ADD_1478 replaced by ADD_5756

//ADD_1477 replaced by ADD_4153

//ADD_1485 replaced by ADD_4223

//ADD_1484 replaced by ADD_5756

//ADD_1483 replaced by ADD_5756

//ADD_1482 replaced by ADD_4158

//ADD_1488 replaced by ADD_4223

//ADD_1487 replaced by ADD_5756

//ADD_1486 replaced by ADD_4162

//ADD_1491 replaced by ADD_4223

//ADD_1490 replaced by ADD_5756

//ADD_1489 replaced by ADD_11602

//ADD_1495 replaced by ADD_4223

//ADD_1494 replaced by ADD_5756

//ADD_1493 replaced by ADD_5756

//ADD_1492 replaced by ADD_4168

//ADD_1499 replaced by ADD_4223

//ADD_1498 replaced by ADD_5756

//ADD_1497 replaced by ADD_5756

//ADD_1496 replaced by ADD_4172

//ADD_1503 replaced by ADD_4223

//ADD_1502 replaced by ADD_5756

//ADD_1501 replaced by ADD_5756

//ADD_1500 replaced by ADD_11602

//ADD_1508 replaced by ADD_4223

//ADD_1507 replaced by ADD_5756

//ADD_1506 replaced by ADD_5756

//ADD_1505 replaced by ADD_5756

//ADD_1504 replaced by ADD_11592

//ADD_1514 replaced by ADD_4223

//ADD_1513 replaced by ADD_5756

//ADD_1512 replaced by ADD_5756

//ADD_1511 replaced by ADD_5756

//ADD_1510 replaced by ADD_5756

//ADD_1509 replaced by ADD_11601

//ADD_1519 replaced by ADD_4223

//ADD_1518 replaced by ADD_5756

//ADD_1517 replaced by ADD_5756

//ADD_1516 replaced by ADD_5756

//ADD_1515 replaced by ADD_4191

//ADD_1524 replaced by ADD_4223

//ADD_1523 replaced by ADD_5756

//ADD_1522 replaced by ADD_5756

//ADD_1521 replaced by ADD_5756

//ADD_1520 replaced by ADD_4196

//ADD_1529 replaced by ADD_4223

//ADD_1528 replaced by ADD_5756

//ADD_1527 replaced by ADD_5756

//ADD_1526 replaced by ADD_5756

//ADD_1525 replaced by ADD_4201

//ADD_1535 replaced by ADD_4223

//ADD_1534 replaced by ADD_5756

//ADD_1533 replaced by ADD_5756

//ADD_1532 replaced by ADD_5756

//ADD_1531 replaced by ADD_5756

//ADD_1530 replaced by ADD_4237

//ADD_1541 replaced by ADD_4223

//ADD_1540 replaced by ADD_5756

//ADD_1539 replaced by ADD_5756

//ADD_1538 replaced by ADD_5756

//ADD_1537 replaced by ADD_5756

//ADD_1536 replaced by ADD_4212

//ADD_1547 replaced by ADD_4223

//ADD_1546 replaced by ADD_5756

//ADD_1545 replaced by ADD_5756

//ADD_1544 replaced by ADD_5756

//ADD_1543 replaced by ADD_5756

//ADD_1542 replaced by ADD_4218

//ADD_1550 replaced by ADD_4226

//ADD_1549 replaced by ADD_5756

//ADD_1548 replaced by ADD_5756

//ADD_1555 replaced by ADD_4231

//ADD_1554 replaced by ADD_5756

//ADD_1553 replaced by ADD_5756

//ADD_1552 replaced by ADD_5756

//ADD_1551 replaced by ADD_5756

//ADD_1561 replaced by ADD_4237

//ADD_1560 replaced by ADD_5756

//ADD_1559 replaced by ADD_5756

//ADD_1558 replaced by ADD_5756

//ADD_1557 replaced by ADD_5756

//ADD_1556 replaced by ADD_5756

//ADD_1567 replaced by ADD_11592

//ADD_1566 replaced by ADD_5756

//ADD_1565 replaced by ADD_5756

//ADD_1564 replaced by ADD_5756

//ADD_1563 replaced by ADD_5756

//ADD_1562 replaced by ADD_5756

//BADD_1225 replaced by BADD_1312

//BADD_1224 replaced by BADD_1311

//BADD_1223 replaced by BADD_1310

//ADD_1575 replaced by ADD_11602

//ADD_1574 replaced by ADD_11602

//ADD_1573 replaced by ADD_11602

//ADD_1572 replaced by ADD_11602

//ADD_1571 replaced by ADD_11602

//ADD_1570 replaced by ADD_11602

//ADD_1569 replaced by ADD_11602

//ADD_1568 replaced by ADD_11602

//KaratsubaCore_68 replaced by KaratsubaCore_143

//KaratsubaCore_67 replaced by KaratsubaCore_142

//KaratsubaCore_66 replaced by KaratsubaCore_141

//BADD_1228 replaced by BADD_1312

//BADD_1227 replaced by BADD_1311

//BADD_1226 replaced by BADD_1310

//ADD_1583 replaced by ADD_11602

//ADD_1582 replaced by ADD_11602

//ADD_1581 replaced by ADD_11602

//ADD_1580 replaced by ADD_11602

//ADD_1579 replaced by ADD_11602

//ADD_1578 replaced by ADD_11602

//ADD_1577 replaced by ADD_11602

//ADD_1576 replaced by ADD_11602

//KaratsubaCore_71 replaced by KaratsubaCore_143

//KaratsubaCore_70 replaced by KaratsubaCore_142

//KaratsubaCore_69 replaced by KaratsubaCore_141

//BADD_1229 replaced by BADD_1306

//ADD_1589 replaced by ADD_5761

//ADD_1588 replaced by ADD_5756

//ADD_1587 replaced by ADD_5756

//ADD_1586 replaced by ADD_5756

//ADD_1585 replaced by ADD_5756

//ADD_1584 replaced by ADD_5756

//ADD_1595 replaced by ADD_4223

//ADD_1594 replaced by ADD_5756

//ADD_1593 replaced by ADD_5756

//ADD_1592 replaced by ADD_5756

//ADD_1591 replaced by ADD_5756

//ADD_1590 replaced by ADD_5756

//ADD_1597 replaced by ADD_4223

//ADD_1596 replaced by ADD_4226

//ADD_1598 replaced by ADD_4055

//ADD_1599 replaced by ADD_4057

//ADD_1601 replaced by ADD_4223

//ADD_1600 replaced by ADD_4057

//ADD_1602 replaced by ADD_4223

//ADD_1603 replaced by ADD_4060

//ADD_1605 replaced by ADD_4223

//ADD_1604 replaced by ADD_11560

//ADD_1607 replaced by ADD_4223

//ADD_1606 replaced by ADD_4196

//ADD_1609 replaced by ADD_4223

//ADD_1608 replaced by ADD_4132

//ADD_1611 replaced by ADD_4223

//ADD_1610 replaced by ADD_4067

//ADD_1615 replaced by ADD_4223

//ADD_1614 replaced by ADD_5756

//ADD_1613 replaced by ADD_5756

//ADD_1612 replaced by ADD_11592

//ADD_1618 replaced by ADD_4223

//ADD_1617 replaced by ADD_5756

//ADD_1616 replaced by ADD_4168

//ADD_1621 replaced by ADD_4223

//ADD_1620 replaced by ADD_5756

//ADD_1619 replaced by ADD_4076

//ADD_1624 replaced by ADD_4223

//ADD_1623 replaced by ADD_5756

//ADD_1622 replaced by ADD_11592

//ADD_1627 replaced by ADD_4223

//ADD_1626 replaced by ADD_5756

//ADD_1625 replaced by ADD_4106

//ADD_1630 replaced by ADD_4223

//ADD_1629 replaced by ADD_5756

//ADD_1628 replaced by ADD_4085

//ADD_1633 replaced by ADD_4223

//ADD_1632 replaced by ADD_5756

//ADD_1631 replaced by ADD_4158

//ADD_1636 replaced by ADD_4223

//ADD_1635 replaced by ADD_5756

//ADD_1634 replaced by ADD_4091

//ADD_1640 replaced by ADD_4223

//ADD_1639 replaced by ADD_5756

//ADD_1638 replaced by ADD_5756

//ADD_1637 replaced by ADD_4094

//ADD_1644 replaced by ADD_4223

//ADD_1643 replaced by ADD_5756

//ADD_1642 replaced by ADD_5756

//ADD_1641 replaced by ADD_4145

//ADD_1648 replaced by ADD_4223

//ADD_1647 replaced by ADD_5756

//ADD_1646 replaced by ADD_5756

//ADD_1645 replaced by ADD_4212

//ADD_1652 replaced by ADD_4223

//ADD_1651 replaced by ADD_5756

//ADD_1650 replaced by ADD_5756

//ADD_1649 replaced by ADD_4106

//ADD_1657 replaced by ADD_4223

//ADD_1656 replaced by ADD_5756

//ADD_1655 replaced by ADD_5756

//ADD_1654 replaced by ADD_5756

//ADD_1653 replaced by ADD_4212

//ADD_1661 replaced by ADD_4223

//ADD_1660 replaced by ADD_5756

//ADD_1659 replaced by ADD_5756

//ADD_1658 replaced by ADD_4115

//ADD_1666 replaced by ADD_4223

//ADD_1665 replaced by ADD_5756

//ADD_1664 replaced by ADD_5756

//ADD_1663 replaced by ADD_5756

//ADD_1662 replaced by ADD_4231

//ADD_1667 replaced by ADD_11560

//ADD_1670 replaced by ADD_4223

//ADD_1669 replaced by ADD_5756

//ADD_1668 replaced by ADD_4125

//ADD_1672 replaced by ADD_4223

//ADD_1671 replaced by ADD_4131

//ADD_1673 replaced by ADD_4150

//ADD_1674 replaced by ADD_4131

//ADD_1675 replaced by ADD_4132

//ADD_1676 replaced by ADD_4196

//ADD_1677 replaced by ADD_4134

//ADD_1678 replaced by ADD_4139

//ADD_1679 replaced by ADD_4136

//ADD_1681 replaced by ADD_4223

//ADD_1680 replaced by ADD_4172

//ADD_1683 replaced by ADD_4223

//ADD_1682 replaced by ADD_4139

//ADD_1685 replaced by ADD_4223

//ADD_1684 replaced by ADD_4141

//ADD_1687 replaced by ADD_4223

//ADD_1686 replaced by ADD_11602

//ADD_1690 replaced by ADD_4223

//ADD_1689 replaced by ADD_5756

//ADD_1688 replaced by ADD_4145

//ADD_1692 replaced by ADD_4223

//ADD_1691 replaced by ADD_5761

//ADD_1695 replaced by ADD_4223

//ADD_1694 replaced by ADD_5756

//ADD_1693 replaced by ADD_4150

//ADD_1700 replaced by ADD_4223

//ADD_1699 replaced by ADD_5756

//ADD_1698 replaced by ADD_5756

//ADD_1697 replaced by ADD_5756

//ADD_1696 replaced by ADD_4153

//ADD_1704 replaced by ADD_4223

//ADD_1703 replaced by ADD_5756

//ADD_1702 replaced by ADD_5756

//ADD_1701 replaced by ADD_4158

//ADD_1707 replaced by ADD_4223

//ADD_1706 replaced by ADD_5756

//ADD_1705 replaced by ADD_4162

//ADD_1710 replaced by ADD_4223

//ADD_1709 replaced by ADD_5756

//ADD_1708 replaced by ADD_11602

//ADD_1714 replaced by ADD_4223

//ADD_1713 replaced by ADD_5756

//ADD_1712 replaced by ADD_5756

//ADD_1711 replaced by ADD_4168

//ADD_1718 replaced by ADD_4223

//ADD_1717 replaced by ADD_5756

//ADD_1716 replaced by ADD_5756

//ADD_1715 replaced by ADD_4172

//ADD_1722 replaced by ADD_4223

//ADD_1721 replaced by ADD_5756

//ADD_1720 replaced by ADD_5756

//ADD_1719 replaced by ADD_11602

//ADD_1727 replaced by ADD_4223

//ADD_1726 replaced by ADD_5756

//ADD_1725 replaced by ADD_5756

//ADD_1724 replaced by ADD_5756

//ADD_1723 replaced by ADD_11592

//ADD_1733 replaced by ADD_4223

//ADD_1732 replaced by ADD_5756

//ADD_1731 replaced by ADD_5756

//ADD_1730 replaced by ADD_5756

//ADD_1729 replaced by ADD_5756

//ADD_1728 replaced by ADD_11601

//ADD_1738 replaced by ADD_4223

//ADD_1737 replaced by ADD_5756

//ADD_1736 replaced by ADD_5756

//ADD_1735 replaced by ADD_5756

//ADD_1734 replaced by ADD_4191

//ADD_1743 replaced by ADD_4223

//ADD_1742 replaced by ADD_5756

//ADD_1741 replaced by ADD_5756

//ADD_1740 replaced by ADD_5756

//ADD_1739 replaced by ADD_4196

//ADD_1748 replaced by ADD_4223

//ADD_1747 replaced by ADD_5756

//ADD_1746 replaced by ADD_5756

//ADD_1745 replaced by ADD_5756

//ADD_1744 replaced by ADD_4201

//ADD_1754 replaced by ADD_4223

//ADD_1753 replaced by ADD_5756

//ADD_1752 replaced by ADD_5756

//ADD_1751 replaced by ADD_5756

//ADD_1750 replaced by ADD_5756

//ADD_1749 replaced by ADD_4237

//ADD_1760 replaced by ADD_4223

//ADD_1759 replaced by ADD_5756

//ADD_1758 replaced by ADD_5756

//ADD_1757 replaced by ADD_5756

//ADD_1756 replaced by ADD_5756

//ADD_1755 replaced by ADD_4212

//ADD_1766 replaced by ADD_4223

//ADD_1765 replaced by ADD_5756

//ADD_1764 replaced by ADD_5756

//ADD_1763 replaced by ADD_5756

//ADD_1762 replaced by ADD_5756

//ADD_1761 replaced by ADD_4218

//ADD_1769 replaced by ADD_4226

//ADD_1768 replaced by ADD_5756

//ADD_1767 replaced by ADD_5756

//ADD_1774 replaced by ADD_4231

//ADD_1773 replaced by ADD_5756

//ADD_1772 replaced by ADD_5756

//ADD_1771 replaced by ADD_5756

//ADD_1770 replaced by ADD_5756

//ADD_1780 replaced by ADD_4237

//ADD_1779 replaced by ADD_5756

//ADD_1778 replaced by ADD_5756

//ADD_1777 replaced by ADD_5756

//ADD_1776 replaced by ADD_5756

//ADD_1775 replaced by ADD_5756

//ADD_1786 replaced by ADD_11592

//ADD_1785 replaced by ADD_5756

//ADD_1784 replaced by ADD_5756

//ADD_1783 replaced by ADD_5756

//ADD_1782 replaced by ADD_5756

//ADD_1781 replaced by ADD_5756

//BADD_1232 replaced by BADD_1312

//BADD_1231 replaced by BADD_1311

//BADD_1230 replaced by BADD_1310

//ADD_1794 replaced by ADD_11602

//ADD_1793 replaced by ADD_11602

//ADD_1792 replaced by ADD_11602

//ADD_1791 replaced by ADD_11602

//ADD_1790 replaced by ADD_11602

//ADD_1789 replaced by ADD_11602

//ADD_1788 replaced by ADD_11602

//ADD_1787 replaced by ADD_11602

//KaratsubaCore_74 replaced by KaratsubaCore_143

//KaratsubaCore_73 replaced by KaratsubaCore_142

//KaratsubaCore_72 replaced by KaratsubaCore_141

//BADD_1235 replaced by BADD_1312

//BADD_1234 replaced by BADD_1311

//BADD_1233 replaced by BADD_1310

//ADD_1802 replaced by ADD_11602

//ADD_1801 replaced by ADD_11602

//ADD_1800 replaced by ADD_11602

//ADD_1799 replaced by ADD_11602

//ADD_1798 replaced by ADD_11602

//ADD_1797 replaced by ADD_11602

//ADD_1796 replaced by ADD_11602

//ADD_1795 replaced by ADD_11602

//KaratsubaCore_77 replaced by KaratsubaCore_143

//KaratsubaCore_76 replaced by KaratsubaCore_142

//KaratsubaCore_75 replaced by KaratsubaCore_141

//BADD_1236 replaced by BADD_1306

//ADD_1808 replaced by ADD_5761

//ADD_1807 replaced by ADD_5756

//ADD_1806 replaced by ADD_5756

//ADD_1805 replaced by ADD_5756

//ADD_1804 replaced by ADD_5756

//ADD_1803 replaced by ADD_5756

//ADD_1814 replaced by ADD_4223

//ADD_1813 replaced by ADD_5756

//ADD_1812 replaced by ADD_5756

//ADD_1811 replaced by ADD_5756

//ADD_1810 replaced by ADD_5756

//ADD_1809 replaced by ADD_5756

//ADD_1816 replaced by ADD_4223

//ADD_1815 replaced by ADD_4226

//ADD_1817 replaced by ADD_4055

//ADD_1818 replaced by ADD_4057

//ADD_1820 replaced by ADD_4223

//ADD_1819 replaced by ADD_4057

//ADD_1821 replaced by ADD_4223

//ADD_1822 replaced by ADD_4060

//ADD_1824 replaced by ADD_4223

//ADD_1823 replaced by ADD_11560

//ADD_1826 replaced by ADD_4223

//ADD_1825 replaced by ADD_4196

//ADD_1828 replaced by ADD_4223

//ADD_1827 replaced by ADD_4132

//ADD_1830 replaced by ADD_4223

//ADD_1829 replaced by ADD_4067

//ADD_1834 replaced by ADD_4223

//ADD_1833 replaced by ADD_5756

//ADD_1832 replaced by ADD_5756

//ADD_1831 replaced by ADD_11592

//ADD_1837 replaced by ADD_4223

//ADD_1836 replaced by ADD_5756

//ADD_1835 replaced by ADD_4168

//ADD_1840 replaced by ADD_4223

//ADD_1839 replaced by ADD_5756

//ADD_1838 replaced by ADD_4076

//ADD_1843 replaced by ADD_4223

//ADD_1842 replaced by ADD_5756

//ADD_1841 replaced by ADD_11592

//ADD_1846 replaced by ADD_4223

//ADD_1845 replaced by ADD_5756

//ADD_1844 replaced by ADD_4106

//ADD_1849 replaced by ADD_4223

//ADD_1848 replaced by ADD_5756

//ADD_1847 replaced by ADD_4085

//ADD_1852 replaced by ADD_4223

//ADD_1851 replaced by ADD_5756

//ADD_1850 replaced by ADD_4158

//ADD_1855 replaced by ADD_4223

//ADD_1854 replaced by ADD_5756

//ADD_1853 replaced by ADD_4091

//ADD_1859 replaced by ADD_4223

//ADD_1858 replaced by ADD_5756

//ADD_1857 replaced by ADD_5756

//ADD_1856 replaced by ADD_4094

//ADD_1863 replaced by ADD_4223

//ADD_1862 replaced by ADD_5756

//ADD_1861 replaced by ADD_5756

//ADD_1860 replaced by ADD_4145

//ADD_1867 replaced by ADD_4223

//ADD_1866 replaced by ADD_5756

//ADD_1865 replaced by ADD_5756

//ADD_1864 replaced by ADD_4212

//ADD_1871 replaced by ADD_4223

//ADD_1870 replaced by ADD_5756

//ADD_1869 replaced by ADD_5756

//ADD_1868 replaced by ADD_4106

//ADD_1876 replaced by ADD_4223

//ADD_1875 replaced by ADD_5756

//ADD_1874 replaced by ADD_5756

//ADD_1873 replaced by ADD_5756

//ADD_1872 replaced by ADD_4212

//ADD_1880 replaced by ADD_4223

//ADD_1879 replaced by ADD_5756

//ADD_1878 replaced by ADD_5756

//ADD_1877 replaced by ADD_4115

//ADD_1885 replaced by ADD_4223

//ADD_1884 replaced by ADD_5756

//ADD_1883 replaced by ADD_5756

//ADD_1882 replaced by ADD_5756

//ADD_1881 replaced by ADD_4231

//ADD_1886 replaced by ADD_11560

//ADD_1889 replaced by ADD_4223

//ADD_1888 replaced by ADD_5756

//ADD_1887 replaced by ADD_4125

//ADD_1891 replaced by ADD_4223

//ADD_1890 replaced by ADD_4131

//ADD_1892 replaced by ADD_4150

//ADD_1893 replaced by ADD_4131

//ADD_1894 replaced by ADD_4132

//ADD_1895 replaced by ADD_4196

//ADD_1896 replaced by ADD_4134

//ADD_1897 replaced by ADD_4139

//ADD_1898 replaced by ADD_4136

//ADD_1900 replaced by ADD_4223

//ADD_1899 replaced by ADD_4172

//ADD_1902 replaced by ADD_4223

//ADD_1901 replaced by ADD_4139

//ADD_1904 replaced by ADD_4223

//ADD_1903 replaced by ADD_4141

//ADD_1906 replaced by ADD_4223

//ADD_1905 replaced by ADD_11602

//ADD_1909 replaced by ADD_4223

//ADD_1908 replaced by ADD_5756

//ADD_1907 replaced by ADD_4145

//ADD_1911 replaced by ADD_4223

//ADD_1910 replaced by ADD_5761

//ADD_1914 replaced by ADD_4223

//ADD_1913 replaced by ADD_5756

//ADD_1912 replaced by ADD_4150

//ADD_1919 replaced by ADD_4223

//ADD_1918 replaced by ADD_5756

//ADD_1917 replaced by ADD_5756

//ADD_1916 replaced by ADD_5756

//ADD_1915 replaced by ADD_4153

//ADD_1923 replaced by ADD_4223

//ADD_1922 replaced by ADD_5756

//ADD_1921 replaced by ADD_5756

//ADD_1920 replaced by ADD_4158

//ADD_1926 replaced by ADD_4223

//ADD_1925 replaced by ADD_5756

//ADD_1924 replaced by ADD_4162

//ADD_1929 replaced by ADD_4223

//ADD_1928 replaced by ADD_5756

//ADD_1927 replaced by ADD_11602

//ADD_1933 replaced by ADD_4223

//ADD_1932 replaced by ADD_5756

//ADD_1931 replaced by ADD_5756

//ADD_1930 replaced by ADD_4168

//ADD_1937 replaced by ADD_4223

//ADD_1936 replaced by ADD_5756

//ADD_1935 replaced by ADD_5756

//ADD_1934 replaced by ADD_4172

//ADD_1941 replaced by ADD_4223

//ADD_1940 replaced by ADD_5756

//ADD_1939 replaced by ADD_5756

//ADD_1938 replaced by ADD_11602

//ADD_1946 replaced by ADD_4223

//ADD_1945 replaced by ADD_5756

//ADD_1944 replaced by ADD_5756

//ADD_1943 replaced by ADD_5756

//ADD_1942 replaced by ADD_11592

//ADD_1952 replaced by ADD_4223

//ADD_1951 replaced by ADD_5756

//ADD_1950 replaced by ADD_5756

//ADD_1949 replaced by ADD_5756

//ADD_1948 replaced by ADD_5756

//ADD_1947 replaced by ADD_11601

//ADD_1957 replaced by ADD_4223

//ADD_1956 replaced by ADD_5756

//ADD_1955 replaced by ADD_5756

//ADD_1954 replaced by ADD_5756

//ADD_1953 replaced by ADD_4191

//ADD_1962 replaced by ADD_4223

//ADD_1961 replaced by ADD_5756

//ADD_1960 replaced by ADD_5756

//ADD_1959 replaced by ADD_5756

//ADD_1958 replaced by ADD_4196

//ADD_1967 replaced by ADD_4223

//ADD_1966 replaced by ADD_5756

//ADD_1965 replaced by ADD_5756

//ADD_1964 replaced by ADD_5756

//ADD_1963 replaced by ADD_4201

//ADD_1973 replaced by ADD_4223

//ADD_1972 replaced by ADD_5756

//ADD_1971 replaced by ADD_5756

//ADD_1970 replaced by ADD_5756

//ADD_1969 replaced by ADD_5756

//ADD_1968 replaced by ADD_4237

//ADD_1979 replaced by ADD_4223

//ADD_1978 replaced by ADD_5756

//ADD_1977 replaced by ADD_5756

//ADD_1976 replaced by ADD_5756

//ADD_1975 replaced by ADD_5756

//ADD_1974 replaced by ADD_4212

//ADD_1985 replaced by ADD_4223

//ADD_1984 replaced by ADD_5756

//ADD_1983 replaced by ADD_5756

//ADD_1982 replaced by ADD_5756

//ADD_1981 replaced by ADD_5756

//ADD_1980 replaced by ADD_4218

//ADD_1988 replaced by ADD_4226

//ADD_1987 replaced by ADD_5756

//ADD_1986 replaced by ADD_5756

//ADD_1993 replaced by ADD_4231

//ADD_1992 replaced by ADD_5756

//ADD_1991 replaced by ADD_5756

//ADD_1990 replaced by ADD_5756

//ADD_1989 replaced by ADD_5756

//ADD_1999 replaced by ADD_4237

//ADD_1998 replaced by ADD_5756

//ADD_1997 replaced by ADD_5756

//ADD_1996 replaced by ADD_5756

//ADD_1995 replaced by ADD_5756

//ADD_1994 replaced by ADD_5756

//ADD_2005 replaced by ADD_11592

//ADD_2004 replaced by ADD_5756

//ADD_2003 replaced by ADD_5756

//ADD_2002 replaced by ADD_5756

//ADD_2001 replaced by ADD_5756

//ADD_2000 replaced by ADD_5756

//BADD_1239 replaced by BADD_1312

//BADD_1238 replaced by BADD_1311

//BADD_1237 replaced by BADD_1310

//ADD_2013 replaced by ADD_11602

//ADD_2012 replaced by ADD_11602

//ADD_2011 replaced by ADD_11602

//ADD_2010 replaced by ADD_11602

//ADD_2009 replaced by ADD_11602

//ADD_2008 replaced by ADD_11602

//ADD_2007 replaced by ADD_11602

//ADD_2006 replaced by ADD_11602

//KaratsubaCore_80 replaced by KaratsubaCore_143

//KaratsubaCore_79 replaced by KaratsubaCore_142

//KaratsubaCore_78 replaced by KaratsubaCore_141

//BADD_1242 replaced by BADD_1312

//BADD_1241 replaced by BADD_1311

//BADD_1240 replaced by BADD_1310

//ADD_2021 replaced by ADD_11602

//ADD_2020 replaced by ADD_11602

//ADD_2019 replaced by ADD_11602

//ADD_2018 replaced by ADD_11602

//ADD_2017 replaced by ADD_11602

//ADD_2016 replaced by ADD_11602

//ADD_2015 replaced by ADD_11602

//ADD_2014 replaced by ADD_11602

//KaratsubaCore_83 replaced by KaratsubaCore_143

//KaratsubaCore_82 replaced by KaratsubaCore_142

//KaratsubaCore_81 replaced by KaratsubaCore_141

//BADD_1243 replaced by BADD_1306

//ADD_2027 replaced by ADD_5761

//ADD_2026 replaced by ADD_5756

//ADD_2025 replaced by ADD_5756

//ADD_2024 replaced by ADD_5756

//ADD_2023 replaced by ADD_5756

//ADD_2022 replaced by ADD_5756

//ADD_2033 replaced by ADD_4223

//ADD_2032 replaced by ADD_5756

//ADD_2031 replaced by ADD_5756

//ADD_2030 replaced by ADD_5756

//ADD_2029 replaced by ADD_5756

//ADD_2028 replaced by ADD_5756

//ADD_2035 replaced by ADD_4223

//ADD_2034 replaced by ADD_4226

//ADD_2036 replaced by ADD_4055

//ADD_2037 replaced by ADD_4057

//ADD_2039 replaced by ADD_4223

//ADD_2038 replaced by ADD_4057

//ADD_2040 replaced by ADD_4223

//ADD_2041 replaced by ADD_4060

//ADD_2043 replaced by ADD_4223

//ADD_2042 replaced by ADD_11560

//ADD_2045 replaced by ADD_4223

//ADD_2044 replaced by ADD_4196

//ADD_2047 replaced by ADD_4223

//ADD_2046 replaced by ADD_4132

//ADD_2049 replaced by ADD_4223

//ADD_2048 replaced by ADD_4067

//ADD_2053 replaced by ADD_4223

//ADD_2052 replaced by ADD_5756

//ADD_2051 replaced by ADD_5756

//ADD_2050 replaced by ADD_11592

//ADD_2056 replaced by ADD_4223

//ADD_2055 replaced by ADD_5756

//ADD_2054 replaced by ADD_4168

//ADD_2059 replaced by ADD_4223

//ADD_2058 replaced by ADD_5756

//ADD_2057 replaced by ADD_4076

//ADD_2062 replaced by ADD_4223

//ADD_2061 replaced by ADD_5756

//ADD_2060 replaced by ADD_11592

//ADD_2065 replaced by ADD_4223

//ADD_2064 replaced by ADD_5756

//ADD_2063 replaced by ADD_4106

//ADD_2068 replaced by ADD_4223

//ADD_2067 replaced by ADD_5756

//ADD_2066 replaced by ADD_4085

//ADD_2071 replaced by ADD_4223

//ADD_2070 replaced by ADD_5756

//ADD_2069 replaced by ADD_4158

//ADD_2074 replaced by ADD_4223

//ADD_2073 replaced by ADD_5756

//ADD_2072 replaced by ADD_4091

//ADD_2078 replaced by ADD_4223

//ADD_2077 replaced by ADD_5756

//ADD_2076 replaced by ADD_5756

//ADD_2075 replaced by ADD_4094

//ADD_2082 replaced by ADD_4223

//ADD_2081 replaced by ADD_5756

//ADD_2080 replaced by ADD_5756

//ADD_2079 replaced by ADD_4145

//ADD_2086 replaced by ADD_4223

//ADD_2085 replaced by ADD_5756

//ADD_2084 replaced by ADD_5756

//ADD_2083 replaced by ADD_4212

//ADD_2090 replaced by ADD_4223

//ADD_2089 replaced by ADD_5756

//ADD_2088 replaced by ADD_5756

//ADD_2087 replaced by ADD_4106

//ADD_2095 replaced by ADD_4223

//ADD_2094 replaced by ADD_5756

//ADD_2093 replaced by ADD_5756

//ADD_2092 replaced by ADD_5756

//ADD_2091 replaced by ADD_4212

//ADD_2099 replaced by ADD_4223

//ADD_2098 replaced by ADD_5756

//ADD_2097 replaced by ADD_5756

//ADD_2096 replaced by ADD_4115

//ADD_2104 replaced by ADD_4223

//ADD_2103 replaced by ADD_5756

//ADD_2102 replaced by ADD_5756

//ADD_2101 replaced by ADD_5756

//ADD_2100 replaced by ADD_4231

//ADD_2105 replaced by ADD_11560

//ADD_2108 replaced by ADD_4223

//ADD_2107 replaced by ADD_5756

//ADD_2106 replaced by ADD_4125

//ADD_2110 replaced by ADD_4223

//ADD_2109 replaced by ADD_4131

//ADD_2111 replaced by ADD_4150

//ADD_2112 replaced by ADD_4131

//ADD_2113 replaced by ADD_4132

//ADD_2114 replaced by ADD_4196

//ADD_2115 replaced by ADD_4134

//ADD_2116 replaced by ADD_4139

//ADD_2117 replaced by ADD_4136

//ADD_2119 replaced by ADD_4223

//ADD_2118 replaced by ADD_4172

//ADD_2121 replaced by ADD_4223

//ADD_2120 replaced by ADD_4139

//ADD_2123 replaced by ADD_4223

//ADD_2122 replaced by ADD_4141

//ADD_2125 replaced by ADD_4223

//ADD_2124 replaced by ADD_11602

//ADD_2128 replaced by ADD_4223

//ADD_2127 replaced by ADD_5756

//ADD_2126 replaced by ADD_4145

//ADD_2130 replaced by ADD_4223

//ADD_2129 replaced by ADD_5761

//ADD_2133 replaced by ADD_4223

//ADD_2132 replaced by ADD_5756

//ADD_2131 replaced by ADD_4150

//ADD_2138 replaced by ADD_4223

//ADD_2137 replaced by ADD_5756

//ADD_2136 replaced by ADD_5756

//ADD_2135 replaced by ADD_5756

//ADD_2134 replaced by ADD_4153

//ADD_2142 replaced by ADD_4223

//ADD_2141 replaced by ADD_5756

//ADD_2140 replaced by ADD_5756

//ADD_2139 replaced by ADD_4158

//ADD_2145 replaced by ADD_4223

//ADD_2144 replaced by ADD_5756

//ADD_2143 replaced by ADD_4162

//ADD_2148 replaced by ADD_4223

//ADD_2147 replaced by ADD_5756

//ADD_2146 replaced by ADD_11602

//ADD_2152 replaced by ADD_4223

//ADD_2151 replaced by ADD_5756

//ADD_2150 replaced by ADD_5756

//ADD_2149 replaced by ADD_4168

//ADD_2156 replaced by ADD_4223

//ADD_2155 replaced by ADD_5756

//ADD_2154 replaced by ADD_5756

//ADD_2153 replaced by ADD_4172

//ADD_2160 replaced by ADD_4223

//ADD_2159 replaced by ADD_5756

//ADD_2158 replaced by ADD_5756

//ADD_2157 replaced by ADD_11602

//ADD_2165 replaced by ADD_4223

//ADD_2164 replaced by ADD_5756

//ADD_2163 replaced by ADD_5756

//ADD_2162 replaced by ADD_5756

//ADD_2161 replaced by ADD_11592

//ADD_2171 replaced by ADD_4223

//ADD_2170 replaced by ADD_5756

//ADD_2169 replaced by ADD_5756

//ADD_2168 replaced by ADD_5756

//ADD_2167 replaced by ADD_5756

//ADD_2166 replaced by ADD_11601

//ADD_2176 replaced by ADD_4223

//ADD_2175 replaced by ADD_5756

//ADD_2174 replaced by ADD_5756

//ADD_2173 replaced by ADD_5756

//ADD_2172 replaced by ADD_4191

//ADD_2181 replaced by ADD_4223

//ADD_2180 replaced by ADD_5756

//ADD_2179 replaced by ADD_5756

//ADD_2178 replaced by ADD_5756

//ADD_2177 replaced by ADD_4196

//ADD_2186 replaced by ADD_4223

//ADD_2185 replaced by ADD_5756

//ADD_2184 replaced by ADD_5756

//ADD_2183 replaced by ADD_5756

//ADD_2182 replaced by ADD_4201

//ADD_2192 replaced by ADD_4223

//ADD_2191 replaced by ADD_5756

//ADD_2190 replaced by ADD_5756

//ADD_2189 replaced by ADD_5756

//ADD_2188 replaced by ADD_5756

//ADD_2187 replaced by ADD_4237

//ADD_2198 replaced by ADD_4223

//ADD_2197 replaced by ADD_5756

//ADD_2196 replaced by ADD_5756

//ADD_2195 replaced by ADD_5756

//ADD_2194 replaced by ADD_5756

//ADD_2193 replaced by ADD_4212

//ADD_2204 replaced by ADD_4223

//ADD_2203 replaced by ADD_5756

//ADD_2202 replaced by ADD_5756

//ADD_2201 replaced by ADD_5756

//ADD_2200 replaced by ADD_5756

//ADD_2199 replaced by ADD_4218

//ADD_2207 replaced by ADD_4226

//ADD_2206 replaced by ADD_5756

//ADD_2205 replaced by ADD_5756

//ADD_2212 replaced by ADD_4231

//ADD_2211 replaced by ADD_5756

//ADD_2210 replaced by ADD_5756

//ADD_2209 replaced by ADD_5756

//ADD_2208 replaced by ADD_5756

//ADD_2218 replaced by ADD_4237

//ADD_2217 replaced by ADD_5756

//ADD_2216 replaced by ADD_5756

//ADD_2215 replaced by ADD_5756

//ADD_2214 replaced by ADD_5756

//ADD_2213 replaced by ADD_5756

//ADD_2224 replaced by ADD_11592

//ADD_2223 replaced by ADD_5756

//ADD_2222 replaced by ADD_5756

//ADD_2221 replaced by ADD_5756

//ADD_2220 replaced by ADD_5756

//ADD_2219 replaced by ADD_5756

//BADD_1246 replaced by BADD_1312

//BADD_1245 replaced by BADD_1311

//BADD_1244 replaced by BADD_1310

//ADD_2232 replaced by ADD_11602

//ADD_2231 replaced by ADD_11602

//ADD_2230 replaced by ADD_11602

//ADD_2229 replaced by ADD_11602

//ADD_2228 replaced by ADD_11602

//ADD_2227 replaced by ADD_11602

//ADD_2226 replaced by ADD_11602

//ADD_2225 replaced by ADD_11602

//KaratsubaCore_86 replaced by KaratsubaCore_143

//KaratsubaCore_85 replaced by KaratsubaCore_142

//KaratsubaCore_84 replaced by KaratsubaCore_141

//BADD_1249 replaced by BADD_1312

//BADD_1248 replaced by BADD_1311

//BADD_1247 replaced by BADD_1310

//ADD_2240 replaced by ADD_11602

//ADD_2239 replaced by ADD_11602

//ADD_2238 replaced by ADD_11602

//ADD_2237 replaced by ADD_11602

//ADD_2236 replaced by ADD_11602

//ADD_2235 replaced by ADD_11602

//ADD_2234 replaced by ADD_11602

//ADD_2233 replaced by ADD_11602

//KaratsubaCore_89 replaced by KaratsubaCore_143

//KaratsubaCore_88 replaced by KaratsubaCore_142

//KaratsubaCore_87 replaced by KaratsubaCore_141

//ADD_2246 replaced by ADD_5761

//ADD_2245 replaced by ADD_5756

//ADD_2244 replaced by ADD_5756

//ADD_2243 replaced by ADD_5756

//ADD_2242 replaced by ADD_5756

//ADD_2241 replaced by ADD_5756

//ADD_2252 replaced by ADD_5761

//ADD_2251 replaced by ADD_5756

//ADD_2250 replaced by ADD_5756

//ADD_2249 replaced by ADD_5756

//ADD_2248 replaced by ADD_5756

//ADD_2247 replaced by ADD_5756

//ADD_2258 replaced by ADD_5761

//ADD_2257 replaced by ADD_5756

//ADD_2256 replaced by ADD_5756

//ADD_2255 replaced by ADD_5756

//ADD_2254 replaced by ADD_5756

//ADD_2253 replaced by ADD_5756

//ADD_2264 replaced by ADD_5761

//ADD_2263 replaced by ADD_5756

//ADD_2262 replaced by ADD_5756

//ADD_2261 replaced by ADD_5756

//ADD_2260 replaced by ADD_5756

//ADD_2259 replaced by ADD_5756

//ADD_2270 replaced by ADD_5761

//ADD_2269 replaced by ADD_5756

//ADD_2268 replaced by ADD_5756

//ADD_2267 replaced by ADD_5756

//ADD_2266 replaced by ADD_5756

//ADD_2265 replaced by ADD_5756

//ADD_2276 replaced by ADD_5761

//ADD_2275 replaced by ADD_5756

//ADD_2274 replaced by ADD_5756

//ADD_2273 replaced by ADD_5756

//ADD_2272 replaced by ADD_5756

//ADD_2271 replaced by ADD_5756

//ADD_2282 replaced by ADD_5761

//ADD_2281 replaced by ADD_5756

//ADD_2280 replaced by ADD_5756

//ADD_2279 replaced by ADD_5756

//ADD_2278 replaced by ADD_5756

//ADD_2277 replaced by ADD_5756

//ADD_2288 replaced by ADD_5761

//ADD_2287 replaced by ADD_5756

//ADD_2286 replaced by ADD_5756

//ADD_2285 replaced by ADD_5756

//ADD_2284 replaced by ADD_5756

//ADD_2283 replaced by ADD_5756

//BADD_1250 replaced by BADD_1306

//ADD_2294 replaced by ADD_5761

//ADD_2293 replaced by ADD_5756

//ADD_2292 replaced by ADD_5756

//ADD_2291 replaced by ADD_5756

//ADD_2290 replaced by ADD_5756

//ADD_2289 replaced by ADD_5756

//ADD_2300 replaced by ADD_4223

//ADD_2299 replaced by ADD_5756

//ADD_2298 replaced by ADD_5756

//ADD_2297 replaced by ADD_5756

//ADD_2296 replaced by ADD_5756

//ADD_2295 replaced by ADD_5756

//ADD_2302 replaced by ADD_4223

//ADD_2301 replaced by ADD_4226

//ADD_2303 replaced by ADD_4055

//ADD_2304 replaced by ADD_4057

//ADD_2306 replaced by ADD_4223

//ADD_2305 replaced by ADD_4057

//ADD_2307 replaced by ADD_4223

//ADD_2308 replaced by ADD_4060

//ADD_2310 replaced by ADD_4223

//ADD_2309 replaced by ADD_11560

//ADD_2312 replaced by ADD_4223

//ADD_2311 replaced by ADD_4196

//ADD_2314 replaced by ADD_4223

//ADD_2313 replaced by ADD_4132

//ADD_2316 replaced by ADD_4223

//ADD_2315 replaced by ADD_4067

//ADD_2320 replaced by ADD_4223

//ADD_2319 replaced by ADD_5756

//ADD_2318 replaced by ADD_5756

//ADD_2317 replaced by ADD_11592

//ADD_2323 replaced by ADD_4223

//ADD_2322 replaced by ADD_5756

//ADD_2321 replaced by ADD_4168

//ADD_2326 replaced by ADD_4223

//ADD_2325 replaced by ADD_5756

//ADD_2324 replaced by ADD_4076

//ADD_2329 replaced by ADD_4223

//ADD_2328 replaced by ADD_5756

//ADD_2327 replaced by ADD_11592

//ADD_2332 replaced by ADD_4223

//ADD_2331 replaced by ADD_5756

//ADD_2330 replaced by ADD_4106

//ADD_2335 replaced by ADD_4223

//ADD_2334 replaced by ADD_5756

//ADD_2333 replaced by ADD_4085

//ADD_2338 replaced by ADD_4223

//ADD_2337 replaced by ADD_5756

//ADD_2336 replaced by ADD_4158

//ADD_2341 replaced by ADD_4223

//ADD_2340 replaced by ADD_5756

//ADD_2339 replaced by ADD_4091

//ADD_2345 replaced by ADD_4223

//ADD_2344 replaced by ADD_5756

//ADD_2343 replaced by ADD_5756

//ADD_2342 replaced by ADD_4094

//ADD_2349 replaced by ADD_4223

//ADD_2348 replaced by ADD_5756

//ADD_2347 replaced by ADD_5756

//ADD_2346 replaced by ADD_4145

//ADD_2353 replaced by ADD_4223

//ADD_2352 replaced by ADD_5756

//ADD_2351 replaced by ADD_5756

//ADD_2350 replaced by ADD_4212

//ADD_2357 replaced by ADD_4223

//ADD_2356 replaced by ADD_5756

//ADD_2355 replaced by ADD_5756

//ADD_2354 replaced by ADD_4106

//ADD_2362 replaced by ADD_4223

//ADD_2361 replaced by ADD_5756

//ADD_2360 replaced by ADD_5756

//ADD_2359 replaced by ADD_5756

//ADD_2358 replaced by ADD_4212

//ADD_2366 replaced by ADD_4223

//ADD_2365 replaced by ADD_5756

//ADD_2364 replaced by ADD_5756

//ADD_2363 replaced by ADD_4115

//ADD_2371 replaced by ADD_4223

//ADD_2370 replaced by ADD_5756

//ADD_2369 replaced by ADD_5756

//ADD_2368 replaced by ADD_5756

//ADD_2367 replaced by ADD_4231

//ADD_2372 replaced by ADD_11560

//ADD_2375 replaced by ADD_4223

//ADD_2374 replaced by ADD_5756

//ADD_2373 replaced by ADD_4125

//ADD_2377 replaced by ADD_4223

//ADD_2376 replaced by ADD_4131

//ADD_2378 replaced by ADD_4150

//ADD_2379 replaced by ADD_4131

//ADD_2380 replaced by ADD_4132

//ADD_2381 replaced by ADD_4196

//ADD_2382 replaced by ADD_4134

//ADD_2383 replaced by ADD_4139

//ADD_2384 replaced by ADD_4136

//ADD_2386 replaced by ADD_4223

//ADD_2385 replaced by ADD_4172

//ADD_2388 replaced by ADD_4223

//ADD_2387 replaced by ADD_4139

//ADD_2390 replaced by ADD_4223

//ADD_2389 replaced by ADD_4141

//ADD_2392 replaced by ADD_4223

//ADD_2391 replaced by ADD_11602

//ADD_2395 replaced by ADD_4223

//ADD_2394 replaced by ADD_5756

//ADD_2393 replaced by ADD_4145

//ADD_2397 replaced by ADD_4223

//ADD_2396 replaced by ADD_5761

//ADD_2400 replaced by ADD_4223

//ADD_2399 replaced by ADD_5756

//ADD_2398 replaced by ADD_4150

//ADD_2405 replaced by ADD_4223

//ADD_2404 replaced by ADD_5756

//ADD_2403 replaced by ADD_5756

//ADD_2402 replaced by ADD_5756

//ADD_2401 replaced by ADD_4153

//ADD_2409 replaced by ADD_4223

//ADD_2408 replaced by ADD_5756

//ADD_2407 replaced by ADD_5756

//ADD_2406 replaced by ADD_4158

//ADD_2412 replaced by ADD_4223

//ADD_2411 replaced by ADD_5756

//ADD_2410 replaced by ADD_4162

//ADD_2415 replaced by ADD_4223

//ADD_2414 replaced by ADD_5756

//ADD_2413 replaced by ADD_11602

//ADD_2419 replaced by ADD_4223

//ADD_2418 replaced by ADD_5756

//ADD_2417 replaced by ADD_5756

//ADD_2416 replaced by ADD_4168

//ADD_2423 replaced by ADD_4223

//ADD_2422 replaced by ADD_5756

//ADD_2421 replaced by ADD_5756

//ADD_2420 replaced by ADD_4172

//ADD_2427 replaced by ADD_4223

//ADD_2426 replaced by ADD_5756

//ADD_2425 replaced by ADD_5756

//ADD_2424 replaced by ADD_11602

//ADD_2432 replaced by ADD_4223

//ADD_2431 replaced by ADD_5756

//ADD_2430 replaced by ADD_5756

//ADD_2429 replaced by ADD_5756

//ADD_2428 replaced by ADD_11592

//ADD_2438 replaced by ADD_4223

//ADD_2437 replaced by ADD_5756

//ADD_2436 replaced by ADD_5756

//ADD_2435 replaced by ADD_5756

//ADD_2434 replaced by ADD_5756

//ADD_2433 replaced by ADD_11601

//ADD_2443 replaced by ADD_4223

//ADD_2442 replaced by ADD_5756

//ADD_2441 replaced by ADD_5756

//ADD_2440 replaced by ADD_5756

//ADD_2439 replaced by ADD_4191

//ADD_2448 replaced by ADD_4223

//ADD_2447 replaced by ADD_5756

//ADD_2446 replaced by ADD_5756

//ADD_2445 replaced by ADD_5756

//ADD_2444 replaced by ADD_4196

//ADD_2453 replaced by ADD_4223

//ADD_2452 replaced by ADD_5756

//ADD_2451 replaced by ADD_5756

//ADD_2450 replaced by ADD_5756

//ADD_2449 replaced by ADD_4201

//ADD_2459 replaced by ADD_4223

//ADD_2458 replaced by ADD_5756

//ADD_2457 replaced by ADD_5756

//ADD_2456 replaced by ADD_5756

//ADD_2455 replaced by ADD_5756

//ADD_2454 replaced by ADD_4237

//ADD_2465 replaced by ADD_4223

//ADD_2464 replaced by ADD_5756

//ADD_2463 replaced by ADD_5756

//ADD_2462 replaced by ADD_5756

//ADD_2461 replaced by ADD_5756

//ADD_2460 replaced by ADD_4212

//ADD_2471 replaced by ADD_4223

//ADD_2470 replaced by ADD_5756

//ADD_2469 replaced by ADD_5756

//ADD_2468 replaced by ADD_5756

//ADD_2467 replaced by ADD_5756

//ADD_2466 replaced by ADD_4218

//ADD_2474 replaced by ADD_4226

//ADD_2473 replaced by ADD_5756

//ADD_2472 replaced by ADD_5756

//ADD_2479 replaced by ADD_4231

//ADD_2478 replaced by ADD_5756

//ADD_2477 replaced by ADD_5756

//ADD_2476 replaced by ADD_5756

//ADD_2475 replaced by ADD_5756

//ADD_2485 replaced by ADD_4237

//ADD_2484 replaced by ADD_5756

//ADD_2483 replaced by ADD_5756

//ADD_2482 replaced by ADD_5756

//ADD_2481 replaced by ADD_5756

//ADD_2480 replaced by ADD_5756

//ADD_2491 replaced by ADD_11592

//ADD_2490 replaced by ADD_5756

//ADD_2489 replaced by ADD_5756

//ADD_2488 replaced by ADD_5756

//ADD_2487 replaced by ADD_5756

//ADD_2486 replaced by ADD_5756

//BADD_1253 replaced by BADD_1312

//BADD_1252 replaced by BADD_1311

//BADD_1251 replaced by BADD_1310

//ADD_2499 replaced by ADD_11602

//ADD_2498 replaced by ADD_11602

//ADD_2497 replaced by ADD_11602

//ADD_2496 replaced by ADD_11602

//ADD_2495 replaced by ADD_11602

//ADD_2494 replaced by ADD_11602

//ADD_2493 replaced by ADD_11602

//ADD_2492 replaced by ADD_11602

//KaratsubaCore_92 replaced by KaratsubaCore_143

//KaratsubaCore_91 replaced by KaratsubaCore_142

//KaratsubaCore_90 replaced by KaratsubaCore_141

//BADD_1256 replaced by BADD_1312

//BADD_1255 replaced by BADD_1311

//BADD_1254 replaced by BADD_1310

//ADD_2507 replaced by ADD_11602

//ADD_2506 replaced by ADD_11602

//ADD_2505 replaced by ADD_11602

//ADD_2504 replaced by ADD_11602

//ADD_2503 replaced by ADD_11602

//ADD_2502 replaced by ADD_11602

//ADD_2501 replaced by ADD_11602

//ADD_2500 replaced by ADD_11602

//KaratsubaCore_95 replaced by KaratsubaCore_143

//KaratsubaCore_94 replaced by KaratsubaCore_142

//KaratsubaCore_93 replaced by KaratsubaCore_141

//BADD_1257 replaced by BADD_1306

//ADD_2513 replaced by ADD_5761

//ADD_2512 replaced by ADD_5756

//ADD_2511 replaced by ADD_5756

//ADD_2510 replaced by ADD_5756

//ADD_2509 replaced by ADD_5756

//ADD_2508 replaced by ADD_5756

//ADD_2519 replaced by ADD_4223

//ADD_2518 replaced by ADD_5756

//ADD_2517 replaced by ADD_5756

//ADD_2516 replaced by ADD_5756

//ADD_2515 replaced by ADD_5756

//ADD_2514 replaced by ADD_5756

//ADD_2521 replaced by ADD_4223

//ADD_2520 replaced by ADD_4226

//ADD_2522 replaced by ADD_4055

//ADD_2523 replaced by ADD_4057

//ADD_2525 replaced by ADD_4223

//ADD_2524 replaced by ADD_4057

//ADD_2526 replaced by ADD_4223

//ADD_2527 replaced by ADD_4060

//ADD_2529 replaced by ADD_4223

//ADD_2528 replaced by ADD_11560

//ADD_2531 replaced by ADD_4223

//ADD_2530 replaced by ADD_4196

//ADD_2533 replaced by ADD_4223

//ADD_2532 replaced by ADD_4132

//ADD_2535 replaced by ADD_4223

//ADD_2534 replaced by ADD_4067

//ADD_2539 replaced by ADD_4223

//ADD_2538 replaced by ADD_5756

//ADD_2537 replaced by ADD_5756

//ADD_2536 replaced by ADD_11592

//ADD_2542 replaced by ADD_4223

//ADD_2541 replaced by ADD_5756

//ADD_2540 replaced by ADD_4168

//ADD_2545 replaced by ADD_4223

//ADD_2544 replaced by ADD_5756

//ADD_2543 replaced by ADD_4076

//ADD_2548 replaced by ADD_4223

//ADD_2547 replaced by ADD_5756

//ADD_2546 replaced by ADD_11592

//ADD_2551 replaced by ADD_4223

//ADD_2550 replaced by ADD_5756

//ADD_2549 replaced by ADD_4106

//ADD_2554 replaced by ADD_4223

//ADD_2553 replaced by ADD_5756

//ADD_2552 replaced by ADD_4085

//ADD_2557 replaced by ADD_4223

//ADD_2556 replaced by ADD_5756

//ADD_2555 replaced by ADD_4158

//ADD_2560 replaced by ADD_4223

//ADD_2559 replaced by ADD_5756

//ADD_2558 replaced by ADD_4091

//ADD_2564 replaced by ADD_4223

//ADD_2563 replaced by ADD_5756

//ADD_2562 replaced by ADD_5756

//ADD_2561 replaced by ADD_4094

//ADD_2568 replaced by ADD_4223

//ADD_2567 replaced by ADD_5756

//ADD_2566 replaced by ADD_5756

//ADD_2565 replaced by ADD_4145

//ADD_2572 replaced by ADD_4223

//ADD_2571 replaced by ADD_5756

//ADD_2570 replaced by ADD_5756

//ADD_2569 replaced by ADD_4212

//ADD_2576 replaced by ADD_4223

//ADD_2575 replaced by ADD_5756

//ADD_2574 replaced by ADD_5756

//ADD_2573 replaced by ADD_4106

//ADD_2581 replaced by ADD_4223

//ADD_2580 replaced by ADD_5756

//ADD_2579 replaced by ADD_5756

//ADD_2578 replaced by ADD_5756

//ADD_2577 replaced by ADD_4212

//ADD_2585 replaced by ADD_4223

//ADD_2584 replaced by ADD_5756

//ADD_2583 replaced by ADD_5756

//ADD_2582 replaced by ADD_4115

//ADD_2590 replaced by ADD_4223

//ADD_2589 replaced by ADD_5756

//ADD_2588 replaced by ADD_5756

//ADD_2587 replaced by ADD_5756

//ADD_2586 replaced by ADD_4231

//ADD_2591 replaced by ADD_11560

//ADD_2594 replaced by ADD_4223

//ADD_2593 replaced by ADD_5756

//ADD_2592 replaced by ADD_4125

//ADD_2596 replaced by ADD_4223

//ADD_2595 replaced by ADD_4131

//ADD_2597 replaced by ADD_4150

//ADD_2598 replaced by ADD_4131

//ADD_2599 replaced by ADD_4132

//ADD_2600 replaced by ADD_4196

//ADD_2601 replaced by ADD_4134

//ADD_2602 replaced by ADD_4139

//ADD_2603 replaced by ADD_4136

//ADD_2605 replaced by ADD_4223

//ADD_2604 replaced by ADD_4172

//ADD_2607 replaced by ADD_4223

//ADD_2606 replaced by ADD_4139

//ADD_2609 replaced by ADD_4223

//ADD_2608 replaced by ADD_4141

//ADD_2611 replaced by ADD_4223

//ADD_2610 replaced by ADD_11602

//ADD_2614 replaced by ADD_4223

//ADD_2613 replaced by ADD_5756

//ADD_2612 replaced by ADD_4145

//ADD_2616 replaced by ADD_4223

//ADD_2615 replaced by ADD_5761

//ADD_2619 replaced by ADD_4223

//ADD_2618 replaced by ADD_5756

//ADD_2617 replaced by ADD_4150

//ADD_2624 replaced by ADD_4223

//ADD_2623 replaced by ADD_5756

//ADD_2622 replaced by ADD_5756

//ADD_2621 replaced by ADD_5756

//ADD_2620 replaced by ADD_4153

//ADD_2628 replaced by ADD_4223

//ADD_2627 replaced by ADD_5756

//ADD_2626 replaced by ADD_5756

//ADD_2625 replaced by ADD_4158

//ADD_2631 replaced by ADD_4223

//ADD_2630 replaced by ADD_5756

//ADD_2629 replaced by ADD_4162

//ADD_2634 replaced by ADD_4223

//ADD_2633 replaced by ADD_5756

//ADD_2632 replaced by ADD_11602

//ADD_2638 replaced by ADD_4223

//ADD_2637 replaced by ADD_5756

//ADD_2636 replaced by ADD_5756

//ADD_2635 replaced by ADD_4168

//ADD_2642 replaced by ADD_4223

//ADD_2641 replaced by ADD_5756

//ADD_2640 replaced by ADD_5756

//ADD_2639 replaced by ADD_4172

//ADD_2646 replaced by ADD_4223

//ADD_2645 replaced by ADD_5756

//ADD_2644 replaced by ADD_5756

//ADD_2643 replaced by ADD_11602

//ADD_2651 replaced by ADD_4223

//ADD_2650 replaced by ADD_5756

//ADD_2649 replaced by ADD_5756

//ADD_2648 replaced by ADD_5756

//ADD_2647 replaced by ADD_11592

//ADD_2657 replaced by ADD_4223

//ADD_2656 replaced by ADD_5756

//ADD_2655 replaced by ADD_5756

//ADD_2654 replaced by ADD_5756

//ADD_2653 replaced by ADD_5756

//ADD_2652 replaced by ADD_11601

//ADD_2662 replaced by ADD_4223

//ADD_2661 replaced by ADD_5756

//ADD_2660 replaced by ADD_5756

//ADD_2659 replaced by ADD_5756

//ADD_2658 replaced by ADD_4191

//ADD_2667 replaced by ADD_4223

//ADD_2666 replaced by ADD_5756

//ADD_2665 replaced by ADD_5756

//ADD_2664 replaced by ADD_5756

//ADD_2663 replaced by ADD_4196

//ADD_2672 replaced by ADD_4223

//ADD_2671 replaced by ADD_5756

//ADD_2670 replaced by ADD_5756

//ADD_2669 replaced by ADD_5756

//ADD_2668 replaced by ADD_4201

//ADD_2678 replaced by ADD_4223

//ADD_2677 replaced by ADD_5756

//ADD_2676 replaced by ADD_5756

//ADD_2675 replaced by ADD_5756

//ADD_2674 replaced by ADD_5756

//ADD_2673 replaced by ADD_4237

//ADD_2684 replaced by ADD_4223

//ADD_2683 replaced by ADD_5756

//ADD_2682 replaced by ADD_5756

//ADD_2681 replaced by ADD_5756

//ADD_2680 replaced by ADD_5756

//ADD_2679 replaced by ADD_4212

//ADD_2690 replaced by ADD_4223

//ADD_2689 replaced by ADD_5756

//ADD_2688 replaced by ADD_5756

//ADD_2687 replaced by ADD_5756

//ADD_2686 replaced by ADD_5756

//ADD_2685 replaced by ADD_4218

//ADD_2693 replaced by ADD_4226

//ADD_2692 replaced by ADD_5756

//ADD_2691 replaced by ADD_5756

//ADD_2698 replaced by ADD_4231

//ADD_2697 replaced by ADD_5756

//ADD_2696 replaced by ADD_5756

//ADD_2695 replaced by ADD_5756

//ADD_2694 replaced by ADD_5756

//ADD_2704 replaced by ADD_4237

//ADD_2703 replaced by ADD_5756

//ADD_2702 replaced by ADD_5756

//ADD_2701 replaced by ADD_5756

//ADD_2700 replaced by ADD_5756

//ADD_2699 replaced by ADD_5756

//ADD_2710 replaced by ADD_11592

//ADD_2709 replaced by ADD_5756

//ADD_2708 replaced by ADD_5756

//ADD_2707 replaced by ADD_5756

//ADD_2706 replaced by ADD_5756

//ADD_2705 replaced by ADD_5756

//BADD_1260 replaced by BADD_1312

//BADD_1259 replaced by BADD_1311

//BADD_1258 replaced by BADD_1310

//ADD_2718 replaced by ADD_11602

//ADD_2717 replaced by ADD_11602

//ADD_2716 replaced by ADD_11602

//ADD_2715 replaced by ADD_11602

//ADD_2714 replaced by ADD_11602

//ADD_2713 replaced by ADD_11602

//ADD_2712 replaced by ADD_11602

//ADD_2711 replaced by ADD_11602

//KaratsubaCore_98 replaced by KaratsubaCore_143

//KaratsubaCore_97 replaced by KaratsubaCore_142

//KaratsubaCore_96 replaced by KaratsubaCore_141

//BADD_1263 replaced by BADD_1312

//BADD_1262 replaced by BADD_1311

//BADD_1261 replaced by BADD_1310

//ADD_2726 replaced by ADD_11602

//ADD_2725 replaced by ADD_11602

//ADD_2724 replaced by ADD_11602

//ADD_2723 replaced by ADD_11602

//ADD_2722 replaced by ADD_11602

//ADD_2721 replaced by ADD_11602

//ADD_2720 replaced by ADD_11602

//ADD_2719 replaced by ADD_11602

//KaratsubaCore_101 replaced by KaratsubaCore_143

//KaratsubaCore_100 replaced by KaratsubaCore_142

//KaratsubaCore_99 replaced by KaratsubaCore_141

//BADD_1264 replaced by BADD_1306

//ADD_2732 replaced by ADD_5761

//ADD_2731 replaced by ADD_5756

//ADD_2730 replaced by ADD_5756

//ADD_2729 replaced by ADD_5756

//ADD_2728 replaced by ADD_5756

//ADD_2727 replaced by ADD_5756

//ADD_2738 replaced by ADD_4223

//ADD_2737 replaced by ADD_5756

//ADD_2736 replaced by ADD_5756

//ADD_2735 replaced by ADD_5756

//ADD_2734 replaced by ADD_5756

//ADD_2733 replaced by ADD_5756

//ADD_2740 replaced by ADD_4223

//ADD_2739 replaced by ADD_4226

//ADD_2741 replaced by ADD_4055

//ADD_2742 replaced by ADD_4057

//ADD_2744 replaced by ADD_4223

//ADD_2743 replaced by ADD_4057

//ADD_2745 replaced by ADD_4223

//ADD_2746 replaced by ADD_4060

//ADD_2748 replaced by ADD_4223

//ADD_2747 replaced by ADD_11560

//ADD_2750 replaced by ADD_4223

//ADD_2749 replaced by ADD_4196

//ADD_2752 replaced by ADD_4223

//ADD_2751 replaced by ADD_4132

//ADD_2754 replaced by ADD_4223

//ADD_2753 replaced by ADD_4067

//ADD_2758 replaced by ADD_4223

//ADD_2757 replaced by ADD_5756

//ADD_2756 replaced by ADD_5756

//ADD_2755 replaced by ADD_11592

//ADD_2761 replaced by ADD_4223

//ADD_2760 replaced by ADD_5756

//ADD_2759 replaced by ADD_4168

//ADD_2764 replaced by ADD_4223

//ADD_2763 replaced by ADD_5756

//ADD_2762 replaced by ADD_4076

//ADD_2767 replaced by ADD_4223

//ADD_2766 replaced by ADD_5756

//ADD_2765 replaced by ADD_11592

//ADD_2770 replaced by ADD_4223

//ADD_2769 replaced by ADD_5756

//ADD_2768 replaced by ADD_4106

//ADD_2773 replaced by ADD_4223

//ADD_2772 replaced by ADD_5756

//ADD_2771 replaced by ADD_4085

//ADD_2776 replaced by ADD_4223

//ADD_2775 replaced by ADD_5756

//ADD_2774 replaced by ADD_4158

//ADD_2779 replaced by ADD_4223

//ADD_2778 replaced by ADD_5756

//ADD_2777 replaced by ADD_4091

//ADD_2783 replaced by ADD_4223

//ADD_2782 replaced by ADD_5756

//ADD_2781 replaced by ADD_5756

//ADD_2780 replaced by ADD_4094

//ADD_2787 replaced by ADD_4223

//ADD_2786 replaced by ADD_5756

//ADD_2785 replaced by ADD_5756

//ADD_2784 replaced by ADD_4145

//ADD_2791 replaced by ADD_4223

//ADD_2790 replaced by ADD_5756

//ADD_2789 replaced by ADD_5756

//ADD_2788 replaced by ADD_4212

//ADD_2795 replaced by ADD_4223

//ADD_2794 replaced by ADD_5756

//ADD_2793 replaced by ADD_5756

//ADD_2792 replaced by ADD_4106

//ADD_2800 replaced by ADD_4223

//ADD_2799 replaced by ADD_5756

//ADD_2798 replaced by ADD_5756

//ADD_2797 replaced by ADD_5756

//ADD_2796 replaced by ADD_4212

//ADD_2804 replaced by ADD_4223

//ADD_2803 replaced by ADD_5756

//ADD_2802 replaced by ADD_5756

//ADD_2801 replaced by ADD_4115

//ADD_2809 replaced by ADD_4223

//ADD_2808 replaced by ADD_5756

//ADD_2807 replaced by ADD_5756

//ADD_2806 replaced by ADD_5756

//ADD_2805 replaced by ADD_4231

//ADD_2810 replaced by ADD_11560

//ADD_2813 replaced by ADD_4223

//ADD_2812 replaced by ADD_5756

//ADD_2811 replaced by ADD_4125

//ADD_2815 replaced by ADD_4223

//ADD_2814 replaced by ADD_4131

//ADD_2816 replaced by ADD_4150

//ADD_2817 replaced by ADD_4131

//ADD_2818 replaced by ADD_4132

//ADD_2819 replaced by ADD_4196

//ADD_2820 replaced by ADD_4134

//ADD_2821 replaced by ADD_4139

//ADD_2822 replaced by ADD_4136

//ADD_2824 replaced by ADD_4223

//ADD_2823 replaced by ADD_4172

//ADD_2826 replaced by ADD_4223

//ADD_2825 replaced by ADD_4139

//ADD_2828 replaced by ADD_4223

//ADD_2827 replaced by ADD_4141

//ADD_2830 replaced by ADD_4223

//ADD_2829 replaced by ADD_11602

//ADD_2833 replaced by ADD_4223

//ADD_2832 replaced by ADD_5756

//ADD_2831 replaced by ADD_4145

//ADD_2835 replaced by ADD_4223

//ADD_2834 replaced by ADD_5761

//ADD_2838 replaced by ADD_4223

//ADD_2837 replaced by ADD_5756

//ADD_2836 replaced by ADD_4150

//ADD_2843 replaced by ADD_4223

//ADD_2842 replaced by ADD_5756

//ADD_2841 replaced by ADD_5756

//ADD_2840 replaced by ADD_5756

//ADD_2839 replaced by ADD_4153

//ADD_2847 replaced by ADD_4223

//ADD_2846 replaced by ADD_5756

//ADD_2845 replaced by ADD_5756

//ADD_2844 replaced by ADD_4158

//ADD_2850 replaced by ADD_4223

//ADD_2849 replaced by ADD_5756

//ADD_2848 replaced by ADD_4162

//ADD_2853 replaced by ADD_4223

//ADD_2852 replaced by ADD_5756

//ADD_2851 replaced by ADD_11602

//ADD_2857 replaced by ADD_4223

//ADD_2856 replaced by ADD_5756

//ADD_2855 replaced by ADD_5756

//ADD_2854 replaced by ADD_4168

//ADD_2861 replaced by ADD_4223

//ADD_2860 replaced by ADD_5756

//ADD_2859 replaced by ADD_5756

//ADD_2858 replaced by ADD_4172

//ADD_2865 replaced by ADD_4223

//ADD_2864 replaced by ADD_5756

//ADD_2863 replaced by ADD_5756

//ADD_2862 replaced by ADD_11602

//ADD_2870 replaced by ADD_4223

//ADD_2869 replaced by ADD_5756

//ADD_2868 replaced by ADD_5756

//ADD_2867 replaced by ADD_5756

//ADD_2866 replaced by ADD_11592

//ADD_2876 replaced by ADD_4223

//ADD_2875 replaced by ADD_5756

//ADD_2874 replaced by ADD_5756

//ADD_2873 replaced by ADD_5756

//ADD_2872 replaced by ADD_5756

//ADD_2871 replaced by ADD_11601

//ADD_2881 replaced by ADD_4223

//ADD_2880 replaced by ADD_5756

//ADD_2879 replaced by ADD_5756

//ADD_2878 replaced by ADD_5756

//ADD_2877 replaced by ADD_4191

//ADD_2886 replaced by ADD_4223

//ADD_2885 replaced by ADD_5756

//ADD_2884 replaced by ADD_5756

//ADD_2883 replaced by ADD_5756

//ADD_2882 replaced by ADD_4196

//ADD_2891 replaced by ADD_4223

//ADD_2890 replaced by ADD_5756

//ADD_2889 replaced by ADD_5756

//ADD_2888 replaced by ADD_5756

//ADD_2887 replaced by ADD_4201

//ADD_2897 replaced by ADD_4223

//ADD_2896 replaced by ADD_5756

//ADD_2895 replaced by ADD_5756

//ADD_2894 replaced by ADD_5756

//ADD_2893 replaced by ADD_5756

//ADD_2892 replaced by ADD_4237

//ADD_2903 replaced by ADD_4223

//ADD_2902 replaced by ADD_5756

//ADD_2901 replaced by ADD_5756

//ADD_2900 replaced by ADD_5756

//ADD_2899 replaced by ADD_5756

//ADD_2898 replaced by ADD_4212

//ADD_2909 replaced by ADD_4223

//ADD_2908 replaced by ADD_5756

//ADD_2907 replaced by ADD_5756

//ADD_2906 replaced by ADD_5756

//ADD_2905 replaced by ADD_5756

//ADD_2904 replaced by ADD_4218

//ADD_2912 replaced by ADD_4226

//ADD_2911 replaced by ADD_5756

//ADD_2910 replaced by ADD_5756

//ADD_2917 replaced by ADD_4231

//ADD_2916 replaced by ADD_5756

//ADD_2915 replaced by ADD_5756

//ADD_2914 replaced by ADD_5756

//ADD_2913 replaced by ADD_5756

//ADD_2923 replaced by ADD_4237

//ADD_2922 replaced by ADD_5756

//ADD_2921 replaced by ADD_5756

//ADD_2920 replaced by ADD_5756

//ADD_2919 replaced by ADD_5756

//ADD_2918 replaced by ADD_5756

//ADD_2929 replaced by ADD_11592

//ADD_2928 replaced by ADD_5756

//ADD_2927 replaced by ADD_5756

//ADD_2926 replaced by ADD_5756

//ADD_2925 replaced by ADD_5756

//ADD_2924 replaced by ADD_5756

//BADD_1267 replaced by BADD_1312

//BADD_1266 replaced by BADD_1311

//BADD_1265 replaced by BADD_1310

//ADD_2937 replaced by ADD_11602

//ADD_2936 replaced by ADD_11602

//ADD_2935 replaced by ADD_11602

//ADD_2934 replaced by ADD_11602

//ADD_2933 replaced by ADD_11602

//ADD_2932 replaced by ADD_11602

//ADD_2931 replaced by ADD_11602

//ADD_2930 replaced by ADD_11602

//KaratsubaCore_104 replaced by KaratsubaCore_143

//KaratsubaCore_103 replaced by KaratsubaCore_142

//KaratsubaCore_102 replaced by KaratsubaCore_141

//BADD_1270 replaced by BADD_1312

//BADD_1269 replaced by BADD_1311

//BADD_1268 replaced by BADD_1310

//ADD_2945 replaced by ADD_11602

//ADD_2944 replaced by ADD_11602

//ADD_2943 replaced by ADD_11602

//ADD_2942 replaced by ADD_11602

//ADD_2941 replaced by ADD_11602

//ADD_2940 replaced by ADD_11602

//ADD_2939 replaced by ADD_11602

//ADD_2938 replaced by ADD_11602

//KaratsubaCore_107 replaced by KaratsubaCore_143

//KaratsubaCore_106 replaced by KaratsubaCore_142

//KaratsubaCore_105 replaced by KaratsubaCore_141

//BADD_1271 replaced by BADD_1306

//ADD_2951 replaced by ADD_5761

//ADD_2950 replaced by ADD_5756

//ADD_2949 replaced by ADD_5756

//ADD_2948 replaced by ADD_5756

//ADD_2947 replaced by ADD_5756

//ADD_2946 replaced by ADD_5756

//ADD_2957 replaced by ADD_4223

//ADD_2956 replaced by ADD_5756

//ADD_2955 replaced by ADD_5756

//ADD_2954 replaced by ADD_5756

//ADD_2953 replaced by ADD_5756

//ADD_2952 replaced by ADD_5756

//ADD_2959 replaced by ADD_4223

//ADD_2958 replaced by ADD_4226

//ADD_2960 replaced by ADD_4055

//ADD_2961 replaced by ADD_4057

//ADD_2963 replaced by ADD_4223

//ADD_2962 replaced by ADD_4057

//ADD_2964 replaced by ADD_4223

//ADD_2965 replaced by ADD_4060

//ADD_2967 replaced by ADD_4223

//ADD_2966 replaced by ADD_11560

//ADD_2969 replaced by ADD_4223

//ADD_2968 replaced by ADD_4196

//ADD_2971 replaced by ADD_4223

//ADD_2970 replaced by ADD_4132

//ADD_2973 replaced by ADD_4223

//ADD_2972 replaced by ADD_4067

//ADD_2977 replaced by ADD_4223

//ADD_2976 replaced by ADD_5756

//ADD_2975 replaced by ADD_5756

//ADD_2974 replaced by ADD_11592

//ADD_2980 replaced by ADD_4223

//ADD_2979 replaced by ADD_5756

//ADD_2978 replaced by ADD_4168

//ADD_2983 replaced by ADD_4223

//ADD_2982 replaced by ADD_5756

//ADD_2981 replaced by ADD_4076

//ADD_2986 replaced by ADD_4223

//ADD_2985 replaced by ADD_5756

//ADD_2984 replaced by ADD_11592

//ADD_2989 replaced by ADD_4223

//ADD_2988 replaced by ADD_5756

//ADD_2987 replaced by ADD_4106

//ADD_2992 replaced by ADD_4223

//ADD_2991 replaced by ADD_5756

//ADD_2990 replaced by ADD_4085

//ADD_2995 replaced by ADD_4223

//ADD_2994 replaced by ADD_5756

//ADD_2993 replaced by ADD_4158

//ADD_2998 replaced by ADD_4223

//ADD_2997 replaced by ADD_5756

//ADD_2996 replaced by ADD_4091

//ADD_3002 replaced by ADD_4223

//ADD_3001 replaced by ADD_5756

//ADD_3000 replaced by ADD_5756

//ADD_2999 replaced by ADD_4094

//ADD_3006 replaced by ADD_4223

//ADD_3005 replaced by ADD_5756

//ADD_3004 replaced by ADD_5756

//ADD_3003 replaced by ADD_4145

//ADD_3010 replaced by ADD_4223

//ADD_3009 replaced by ADD_5756

//ADD_3008 replaced by ADD_5756

//ADD_3007 replaced by ADD_4212

//ADD_3014 replaced by ADD_4223

//ADD_3013 replaced by ADD_5756

//ADD_3012 replaced by ADD_5756

//ADD_3011 replaced by ADD_4106

//ADD_3019 replaced by ADD_4223

//ADD_3018 replaced by ADD_5756

//ADD_3017 replaced by ADD_5756

//ADD_3016 replaced by ADD_5756

//ADD_3015 replaced by ADD_4212

//ADD_3023 replaced by ADD_4223

//ADD_3022 replaced by ADD_5756

//ADD_3021 replaced by ADD_5756

//ADD_3020 replaced by ADD_4115

//ADD_3028 replaced by ADD_4223

//ADD_3027 replaced by ADD_5756

//ADD_3026 replaced by ADD_5756

//ADD_3025 replaced by ADD_5756

//ADD_3024 replaced by ADD_4231

//ADD_3029 replaced by ADD_11560

//ADD_3032 replaced by ADD_4223

//ADD_3031 replaced by ADD_5756

//ADD_3030 replaced by ADD_4125

//ADD_3034 replaced by ADD_4223

//ADD_3033 replaced by ADD_4131

//ADD_3035 replaced by ADD_4150

//ADD_3036 replaced by ADD_4131

//ADD_3037 replaced by ADD_4132

//ADD_3038 replaced by ADD_4196

//ADD_3039 replaced by ADD_4134

//ADD_3040 replaced by ADD_4139

//ADD_3041 replaced by ADD_4136

//ADD_3043 replaced by ADD_4223

//ADD_3042 replaced by ADD_4172

//ADD_3045 replaced by ADD_4223

//ADD_3044 replaced by ADD_4139

//ADD_3047 replaced by ADD_4223

//ADD_3046 replaced by ADD_4141

//ADD_3049 replaced by ADD_4223

//ADD_3048 replaced by ADD_11602

//ADD_3052 replaced by ADD_4223

//ADD_3051 replaced by ADD_5756

//ADD_3050 replaced by ADD_4145

//ADD_3054 replaced by ADD_4223

//ADD_3053 replaced by ADD_5761

//ADD_3057 replaced by ADD_4223

//ADD_3056 replaced by ADD_5756

//ADD_3055 replaced by ADD_4150

//ADD_3062 replaced by ADD_4223

//ADD_3061 replaced by ADD_5756

//ADD_3060 replaced by ADD_5756

//ADD_3059 replaced by ADD_5756

//ADD_3058 replaced by ADD_4153

//ADD_3066 replaced by ADD_4223

//ADD_3065 replaced by ADD_5756

//ADD_3064 replaced by ADD_5756

//ADD_3063 replaced by ADD_4158

//ADD_3069 replaced by ADD_4223

//ADD_3068 replaced by ADD_5756

//ADD_3067 replaced by ADD_4162

//ADD_3072 replaced by ADD_4223

//ADD_3071 replaced by ADD_5756

//ADD_3070 replaced by ADD_11602

//ADD_3076 replaced by ADD_4223

//ADD_3075 replaced by ADD_5756

//ADD_3074 replaced by ADD_5756

//ADD_3073 replaced by ADD_4168

//ADD_3080 replaced by ADD_4223

//ADD_3079 replaced by ADD_5756

//ADD_3078 replaced by ADD_5756

//ADD_3077 replaced by ADD_4172

//ADD_3084 replaced by ADD_4223

//ADD_3083 replaced by ADD_5756

//ADD_3082 replaced by ADD_5756

//ADD_3081 replaced by ADD_11602

//ADD_3089 replaced by ADD_4223

//ADD_3088 replaced by ADD_5756

//ADD_3087 replaced by ADD_5756

//ADD_3086 replaced by ADD_5756

//ADD_3085 replaced by ADD_11592

//ADD_3095 replaced by ADD_4223

//ADD_3094 replaced by ADD_5756

//ADD_3093 replaced by ADD_5756

//ADD_3092 replaced by ADD_5756

//ADD_3091 replaced by ADD_5756

//ADD_3090 replaced by ADD_11601

//ADD_3100 replaced by ADD_4223

//ADD_3099 replaced by ADD_5756

//ADD_3098 replaced by ADD_5756

//ADD_3097 replaced by ADD_5756

//ADD_3096 replaced by ADD_4191

//ADD_3105 replaced by ADD_4223

//ADD_3104 replaced by ADD_5756

//ADD_3103 replaced by ADD_5756

//ADD_3102 replaced by ADD_5756

//ADD_3101 replaced by ADD_4196

//ADD_3110 replaced by ADD_4223

//ADD_3109 replaced by ADD_5756

//ADD_3108 replaced by ADD_5756

//ADD_3107 replaced by ADD_5756

//ADD_3106 replaced by ADD_4201

//ADD_3116 replaced by ADD_4223

//ADD_3115 replaced by ADD_5756

//ADD_3114 replaced by ADD_5756

//ADD_3113 replaced by ADD_5756

//ADD_3112 replaced by ADD_5756

//ADD_3111 replaced by ADD_4237

//ADD_3122 replaced by ADD_4223

//ADD_3121 replaced by ADD_5756

//ADD_3120 replaced by ADD_5756

//ADD_3119 replaced by ADD_5756

//ADD_3118 replaced by ADD_5756

//ADD_3117 replaced by ADD_4212

//ADD_3128 replaced by ADD_4223

//ADD_3127 replaced by ADD_5756

//ADD_3126 replaced by ADD_5756

//ADD_3125 replaced by ADD_5756

//ADD_3124 replaced by ADD_5756

//ADD_3123 replaced by ADD_4218

//ADD_3131 replaced by ADD_4226

//ADD_3130 replaced by ADD_5756

//ADD_3129 replaced by ADD_5756

//ADD_3136 replaced by ADD_4231

//ADD_3135 replaced by ADD_5756

//ADD_3134 replaced by ADD_5756

//ADD_3133 replaced by ADD_5756

//ADD_3132 replaced by ADD_5756

//ADD_3142 replaced by ADD_4237

//ADD_3141 replaced by ADD_5756

//ADD_3140 replaced by ADD_5756

//ADD_3139 replaced by ADD_5756

//ADD_3138 replaced by ADD_5756

//ADD_3137 replaced by ADD_5756

//ADD_3148 replaced by ADD_11592

//ADD_3147 replaced by ADD_5756

//ADD_3146 replaced by ADD_5756

//ADD_3145 replaced by ADD_5756

//ADD_3144 replaced by ADD_5756

//ADD_3143 replaced by ADD_5756

//BADD_1274 replaced by BADD_1312

//BADD_1273 replaced by BADD_1311

//BADD_1272 replaced by BADD_1310

//ADD_3156 replaced by ADD_11602

//ADD_3155 replaced by ADD_11602

//ADD_3154 replaced by ADD_11602

//ADD_3153 replaced by ADD_11602

//ADD_3152 replaced by ADD_11602

//ADD_3151 replaced by ADD_11602

//ADD_3150 replaced by ADD_11602

//ADD_3149 replaced by ADD_11602

//KaratsubaCore_110 replaced by KaratsubaCore_143

//KaratsubaCore_109 replaced by KaratsubaCore_142

//KaratsubaCore_108 replaced by KaratsubaCore_141

//BADD_1277 replaced by BADD_1312

//BADD_1276 replaced by BADD_1311

//BADD_1275 replaced by BADD_1310

//ADD_3164 replaced by ADD_11602

//ADD_3163 replaced by ADD_11602

//ADD_3162 replaced by ADD_11602

//ADD_3161 replaced by ADD_11602

//ADD_3160 replaced by ADD_11602

//ADD_3159 replaced by ADD_11602

//ADD_3158 replaced by ADD_11602

//ADD_3157 replaced by ADD_11602

//KaratsubaCore_113 replaced by KaratsubaCore_143

//KaratsubaCore_112 replaced by KaratsubaCore_142

//KaratsubaCore_111 replaced by KaratsubaCore_141

//BADD_1278 replaced by BADD_1306

//ADD_3170 replaced by ADD_5761

//ADD_3169 replaced by ADD_5756

//ADD_3168 replaced by ADD_5756

//ADD_3167 replaced by ADD_5756

//ADD_3166 replaced by ADD_5756

//ADD_3165 replaced by ADD_5756

//ADD_3176 replaced by ADD_4223

//ADD_3175 replaced by ADD_5756

//ADD_3174 replaced by ADD_5756

//ADD_3173 replaced by ADD_5756

//ADD_3172 replaced by ADD_5756

//ADD_3171 replaced by ADD_5756

//ADD_3178 replaced by ADD_4223

//ADD_3177 replaced by ADD_4226

//ADD_3179 replaced by ADD_4055

//ADD_3180 replaced by ADD_4057

//ADD_3182 replaced by ADD_4223

//ADD_3181 replaced by ADD_4057

//ADD_3183 replaced by ADD_4223

//ADD_3184 replaced by ADD_4060

//ADD_3186 replaced by ADD_4223

//ADD_3185 replaced by ADD_11560

//ADD_3188 replaced by ADD_4223

//ADD_3187 replaced by ADD_4196

//ADD_3190 replaced by ADD_4223

//ADD_3189 replaced by ADD_4132

//ADD_3192 replaced by ADD_4223

//ADD_3191 replaced by ADD_4067

//ADD_3196 replaced by ADD_4223

//ADD_3195 replaced by ADD_5756

//ADD_3194 replaced by ADD_5756

//ADD_3193 replaced by ADD_11592

//ADD_3199 replaced by ADD_4223

//ADD_3198 replaced by ADD_5756

//ADD_3197 replaced by ADD_4168

//ADD_3202 replaced by ADD_4223

//ADD_3201 replaced by ADD_5756

//ADD_3200 replaced by ADD_4076

//ADD_3205 replaced by ADD_4223

//ADD_3204 replaced by ADD_5756

//ADD_3203 replaced by ADD_11592

//ADD_3208 replaced by ADD_4223

//ADD_3207 replaced by ADD_5756

//ADD_3206 replaced by ADD_4106

//ADD_3211 replaced by ADD_4223

//ADD_3210 replaced by ADD_5756

//ADD_3209 replaced by ADD_4085

//ADD_3214 replaced by ADD_4223

//ADD_3213 replaced by ADD_5756

//ADD_3212 replaced by ADD_4158

//ADD_3217 replaced by ADD_4223

//ADD_3216 replaced by ADD_5756

//ADD_3215 replaced by ADD_4091

//ADD_3221 replaced by ADD_4223

//ADD_3220 replaced by ADD_5756

//ADD_3219 replaced by ADD_5756

//ADD_3218 replaced by ADD_4094

//ADD_3225 replaced by ADD_4223

//ADD_3224 replaced by ADD_5756

//ADD_3223 replaced by ADD_5756

//ADD_3222 replaced by ADD_4145

//ADD_3229 replaced by ADD_4223

//ADD_3228 replaced by ADD_5756

//ADD_3227 replaced by ADD_5756

//ADD_3226 replaced by ADD_4212

//ADD_3233 replaced by ADD_4223

//ADD_3232 replaced by ADD_5756

//ADD_3231 replaced by ADD_5756

//ADD_3230 replaced by ADD_4106

//ADD_3238 replaced by ADD_4223

//ADD_3237 replaced by ADD_5756

//ADD_3236 replaced by ADD_5756

//ADD_3235 replaced by ADD_5756

//ADD_3234 replaced by ADD_4212

//ADD_3242 replaced by ADD_4223

//ADD_3241 replaced by ADD_5756

//ADD_3240 replaced by ADD_5756

//ADD_3239 replaced by ADD_4115

//ADD_3247 replaced by ADD_4223

//ADD_3246 replaced by ADD_5756

//ADD_3245 replaced by ADD_5756

//ADD_3244 replaced by ADD_5756

//ADD_3243 replaced by ADD_4231

//ADD_3248 replaced by ADD_11560

//ADD_3251 replaced by ADD_4223

//ADD_3250 replaced by ADD_5756

//ADD_3249 replaced by ADD_4125

//ADD_3253 replaced by ADD_4223

//ADD_3252 replaced by ADD_4131

//ADD_3254 replaced by ADD_4150

//ADD_3255 replaced by ADD_4131

//ADD_3256 replaced by ADD_4132

//ADD_3257 replaced by ADD_4196

//ADD_3258 replaced by ADD_4134

//ADD_3259 replaced by ADD_4139

//ADD_3260 replaced by ADD_4136

//ADD_3262 replaced by ADD_4223

//ADD_3261 replaced by ADD_4172

//ADD_3264 replaced by ADD_4223

//ADD_3263 replaced by ADD_4139

//ADD_3266 replaced by ADD_4223

//ADD_3265 replaced by ADD_4141

//ADD_3268 replaced by ADD_4223

//ADD_3267 replaced by ADD_11602

//ADD_3271 replaced by ADD_4223

//ADD_3270 replaced by ADD_5756

//ADD_3269 replaced by ADD_4145

//ADD_3273 replaced by ADD_4223

//ADD_3272 replaced by ADD_5761

//ADD_3276 replaced by ADD_4223

//ADD_3275 replaced by ADD_5756

//ADD_3274 replaced by ADD_4150

//ADD_3281 replaced by ADD_4223

//ADD_3280 replaced by ADD_5756

//ADD_3279 replaced by ADD_5756

//ADD_3278 replaced by ADD_5756

//ADD_3277 replaced by ADD_4153

//ADD_3285 replaced by ADD_4223

//ADD_3284 replaced by ADD_5756

//ADD_3283 replaced by ADD_5756

//ADD_3282 replaced by ADD_4158

//ADD_3288 replaced by ADD_4223

//ADD_3287 replaced by ADD_5756

//ADD_3286 replaced by ADD_4162

//ADD_3291 replaced by ADD_4223

//ADD_3290 replaced by ADD_5756

//ADD_3289 replaced by ADD_11602

//ADD_3295 replaced by ADD_4223

//ADD_3294 replaced by ADD_5756

//ADD_3293 replaced by ADD_5756

//ADD_3292 replaced by ADD_4168

//ADD_3299 replaced by ADD_4223

//ADD_3298 replaced by ADD_5756

//ADD_3297 replaced by ADD_5756

//ADD_3296 replaced by ADD_4172

//ADD_3303 replaced by ADD_4223

//ADD_3302 replaced by ADD_5756

//ADD_3301 replaced by ADD_5756

//ADD_3300 replaced by ADD_11602

//ADD_3308 replaced by ADD_4223

//ADD_3307 replaced by ADD_5756

//ADD_3306 replaced by ADD_5756

//ADD_3305 replaced by ADD_5756

//ADD_3304 replaced by ADD_11592

//ADD_3314 replaced by ADD_4223

//ADD_3313 replaced by ADD_5756

//ADD_3312 replaced by ADD_5756

//ADD_3311 replaced by ADD_5756

//ADD_3310 replaced by ADD_5756

//ADD_3309 replaced by ADD_11601

//ADD_3319 replaced by ADD_4223

//ADD_3318 replaced by ADD_5756

//ADD_3317 replaced by ADD_5756

//ADD_3316 replaced by ADD_5756

//ADD_3315 replaced by ADD_4191

//ADD_3324 replaced by ADD_4223

//ADD_3323 replaced by ADD_5756

//ADD_3322 replaced by ADD_5756

//ADD_3321 replaced by ADD_5756

//ADD_3320 replaced by ADD_4196

//ADD_3329 replaced by ADD_4223

//ADD_3328 replaced by ADD_5756

//ADD_3327 replaced by ADD_5756

//ADD_3326 replaced by ADD_5756

//ADD_3325 replaced by ADD_4201

//ADD_3335 replaced by ADD_4223

//ADD_3334 replaced by ADD_5756

//ADD_3333 replaced by ADD_5756

//ADD_3332 replaced by ADD_5756

//ADD_3331 replaced by ADD_5756

//ADD_3330 replaced by ADD_4237

//ADD_3341 replaced by ADD_4223

//ADD_3340 replaced by ADD_5756

//ADD_3339 replaced by ADD_5756

//ADD_3338 replaced by ADD_5756

//ADD_3337 replaced by ADD_5756

//ADD_3336 replaced by ADD_4212

//ADD_3347 replaced by ADD_4223

//ADD_3346 replaced by ADD_5756

//ADD_3345 replaced by ADD_5756

//ADD_3344 replaced by ADD_5756

//ADD_3343 replaced by ADD_5756

//ADD_3342 replaced by ADD_4218

//ADD_3350 replaced by ADD_4226

//ADD_3349 replaced by ADD_5756

//ADD_3348 replaced by ADD_5756

//ADD_3355 replaced by ADD_4231

//ADD_3354 replaced by ADD_5756

//ADD_3353 replaced by ADD_5756

//ADD_3352 replaced by ADD_5756

//ADD_3351 replaced by ADD_5756

//ADD_3361 replaced by ADD_4237

//ADD_3360 replaced by ADD_5756

//ADD_3359 replaced by ADD_5756

//ADD_3358 replaced by ADD_5756

//ADD_3357 replaced by ADD_5756

//ADD_3356 replaced by ADD_5756

//ADD_3367 replaced by ADD_11592

//ADD_3366 replaced by ADD_5756

//ADD_3365 replaced by ADD_5756

//ADD_3364 replaced by ADD_5756

//ADD_3363 replaced by ADD_5756

//ADD_3362 replaced by ADD_5756

//BADD_1281 replaced by BADD_1312

//BADD_1280 replaced by BADD_1311

//BADD_1279 replaced by BADD_1310

//ADD_3375 replaced by ADD_11602

//ADD_3374 replaced by ADD_11602

//ADD_3373 replaced by ADD_11602

//ADD_3372 replaced by ADD_11602

//ADD_3371 replaced by ADD_11602

//ADD_3370 replaced by ADD_11602

//ADD_3369 replaced by ADD_11602

//ADD_3368 replaced by ADD_11602

//KaratsubaCore_116 replaced by KaratsubaCore_143

//KaratsubaCore_115 replaced by KaratsubaCore_142

//KaratsubaCore_114 replaced by KaratsubaCore_141

//BADD_1284 replaced by BADD_1312

//BADD_1283 replaced by BADD_1311

//BADD_1282 replaced by BADD_1310

//ADD_3383 replaced by ADD_11602

//ADD_3382 replaced by ADD_11602

//ADD_3381 replaced by ADD_11602

//ADD_3380 replaced by ADD_11602

//ADD_3379 replaced by ADD_11602

//ADD_3378 replaced by ADD_11602

//ADD_3377 replaced by ADD_11602

//ADD_3376 replaced by ADD_11602

//KaratsubaCore_119 replaced by KaratsubaCore_143

//KaratsubaCore_118 replaced by KaratsubaCore_142

//KaratsubaCore_117 replaced by KaratsubaCore_141

//BADD_1285 replaced by BADD_1306

//ADD_3389 replaced by ADD_5761

//ADD_3388 replaced by ADD_5756

//ADD_3387 replaced by ADD_5756

//ADD_3386 replaced by ADD_5756

//ADD_3385 replaced by ADD_5756

//ADD_3384 replaced by ADD_5756

//ADD_3395 replaced by ADD_4223

//ADD_3394 replaced by ADD_5756

//ADD_3393 replaced by ADD_5756

//ADD_3392 replaced by ADD_5756

//ADD_3391 replaced by ADD_5756

//ADD_3390 replaced by ADD_5756

//ADD_3397 replaced by ADD_4223

//ADD_3396 replaced by ADD_4226

//ADD_3398 replaced by ADD_4055

//ADD_3399 replaced by ADD_4057

//ADD_3401 replaced by ADD_4223

//ADD_3400 replaced by ADD_4057

//ADD_3402 replaced by ADD_4223

//ADD_3403 replaced by ADD_4060

//ADD_3405 replaced by ADD_4223

//ADD_3404 replaced by ADD_11560

//ADD_3407 replaced by ADD_4223

//ADD_3406 replaced by ADD_4196

//ADD_3409 replaced by ADD_4223

//ADD_3408 replaced by ADD_4132

//ADD_3411 replaced by ADD_4223

//ADD_3410 replaced by ADD_4067

//ADD_3415 replaced by ADD_4223

//ADD_3414 replaced by ADD_5756

//ADD_3413 replaced by ADD_5756

//ADD_3412 replaced by ADD_11592

//ADD_3418 replaced by ADD_4223

//ADD_3417 replaced by ADD_5756

//ADD_3416 replaced by ADD_4168

//ADD_3421 replaced by ADD_4223

//ADD_3420 replaced by ADD_5756

//ADD_3419 replaced by ADD_4076

//ADD_3424 replaced by ADD_4223

//ADD_3423 replaced by ADD_5756

//ADD_3422 replaced by ADD_11592

//ADD_3427 replaced by ADD_4223

//ADD_3426 replaced by ADD_5756

//ADD_3425 replaced by ADD_4106

//ADD_3430 replaced by ADD_4223

//ADD_3429 replaced by ADD_5756

//ADD_3428 replaced by ADD_4085

//ADD_3433 replaced by ADD_4223

//ADD_3432 replaced by ADD_5756

//ADD_3431 replaced by ADD_4158

//ADD_3436 replaced by ADD_4223

//ADD_3435 replaced by ADD_5756

//ADD_3434 replaced by ADD_4091

//ADD_3440 replaced by ADD_4223

//ADD_3439 replaced by ADD_5756

//ADD_3438 replaced by ADD_5756

//ADD_3437 replaced by ADD_4094

//ADD_3444 replaced by ADD_4223

//ADD_3443 replaced by ADD_5756

//ADD_3442 replaced by ADD_5756

//ADD_3441 replaced by ADD_4145

//ADD_3448 replaced by ADD_4223

//ADD_3447 replaced by ADD_5756

//ADD_3446 replaced by ADD_5756

//ADD_3445 replaced by ADD_4212

//ADD_3452 replaced by ADD_4223

//ADD_3451 replaced by ADD_5756

//ADD_3450 replaced by ADD_5756

//ADD_3449 replaced by ADD_4106

//ADD_3457 replaced by ADD_4223

//ADD_3456 replaced by ADD_5756

//ADD_3455 replaced by ADD_5756

//ADD_3454 replaced by ADD_5756

//ADD_3453 replaced by ADD_4212

//ADD_3461 replaced by ADD_4223

//ADD_3460 replaced by ADD_5756

//ADD_3459 replaced by ADD_5756

//ADD_3458 replaced by ADD_4115

//ADD_3466 replaced by ADD_4223

//ADD_3465 replaced by ADD_5756

//ADD_3464 replaced by ADD_5756

//ADD_3463 replaced by ADD_5756

//ADD_3462 replaced by ADD_4231

//ADD_3467 replaced by ADD_11560

//ADD_3470 replaced by ADD_4223

//ADD_3469 replaced by ADD_5756

//ADD_3468 replaced by ADD_4125

//ADD_3472 replaced by ADD_4223

//ADD_3471 replaced by ADD_4131

//ADD_3473 replaced by ADD_4150

//ADD_3474 replaced by ADD_4131

//ADD_3475 replaced by ADD_4132

//ADD_3476 replaced by ADD_4196

//ADD_3477 replaced by ADD_4134

//ADD_3478 replaced by ADD_4139

//ADD_3479 replaced by ADD_4136

//ADD_3481 replaced by ADD_4223

//ADD_3480 replaced by ADD_4172

//ADD_3483 replaced by ADD_4223

//ADD_3482 replaced by ADD_4139

//ADD_3485 replaced by ADD_4223

//ADD_3484 replaced by ADD_4141

//ADD_3487 replaced by ADD_4223

//ADD_3486 replaced by ADD_11602

//ADD_3490 replaced by ADD_4223

//ADD_3489 replaced by ADD_5756

//ADD_3488 replaced by ADD_4145

//ADD_3492 replaced by ADD_4223

//ADD_3491 replaced by ADD_5761

//ADD_3495 replaced by ADD_4223

//ADD_3494 replaced by ADD_5756

//ADD_3493 replaced by ADD_4150

//ADD_3500 replaced by ADD_4223

//ADD_3499 replaced by ADD_5756

//ADD_3498 replaced by ADD_5756

//ADD_3497 replaced by ADD_5756

//ADD_3496 replaced by ADD_4153

//ADD_3504 replaced by ADD_4223

//ADD_3503 replaced by ADD_5756

//ADD_3502 replaced by ADD_5756

//ADD_3501 replaced by ADD_4158

//ADD_3507 replaced by ADD_4223

//ADD_3506 replaced by ADD_5756

//ADD_3505 replaced by ADD_4162

//ADD_3510 replaced by ADD_4223

//ADD_3509 replaced by ADD_5756

//ADD_3508 replaced by ADD_11602

//ADD_3514 replaced by ADD_4223

//ADD_3513 replaced by ADD_5756

//ADD_3512 replaced by ADD_5756

//ADD_3511 replaced by ADD_4168

//ADD_3518 replaced by ADD_4223

//ADD_3517 replaced by ADD_5756

//ADD_3516 replaced by ADD_5756

//ADD_3515 replaced by ADD_4172

//ADD_3522 replaced by ADD_4223

//ADD_3521 replaced by ADD_5756

//ADD_3520 replaced by ADD_5756

//ADD_3519 replaced by ADD_11602

//ADD_3527 replaced by ADD_4223

//ADD_3526 replaced by ADD_5756

//ADD_3525 replaced by ADD_5756

//ADD_3524 replaced by ADD_5756

//ADD_3523 replaced by ADD_11592

//ADD_3533 replaced by ADD_4223

//ADD_3532 replaced by ADD_5756

//ADD_3531 replaced by ADD_5756

//ADD_3530 replaced by ADD_5756

//ADD_3529 replaced by ADD_5756

//ADD_3528 replaced by ADD_11601

//ADD_3538 replaced by ADD_4223

//ADD_3537 replaced by ADD_5756

//ADD_3536 replaced by ADD_5756

//ADD_3535 replaced by ADD_5756

//ADD_3534 replaced by ADD_4191

//ADD_3543 replaced by ADD_4223

//ADD_3542 replaced by ADD_5756

//ADD_3541 replaced by ADD_5756

//ADD_3540 replaced by ADD_5756

//ADD_3539 replaced by ADD_4196

//ADD_3548 replaced by ADD_4223

//ADD_3547 replaced by ADD_5756

//ADD_3546 replaced by ADD_5756

//ADD_3545 replaced by ADD_5756

//ADD_3544 replaced by ADD_4201

//ADD_3554 replaced by ADD_4223

//ADD_3553 replaced by ADD_5756

//ADD_3552 replaced by ADD_5756

//ADD_3551 replaced by ADD_5756

//ADD_3550 replaced by ADD_5756

//ADD_3549 replaced by ADD_4237

//ADD_3560 replaced by ADD_4223

//ADD_3559 replaced by ADD_5756

//ADD_3558 replaced by ADD_5756

//ADD_3557 replaced by ADD_5756

//ADD_3556 replaced by ADD_5756

//ADD_3555 replaced by ADD_4212

//ADD_3566 replaced by ADD_4223

//ADD_3565 replaced by ADD_5756

//ADD_3564 replaced by ADD_5756

//ADD_3563 replaced by ADD_5756

//ADD_3562 replaced by ADD_5756

//ADD_3561 replaced by ADD_4218

//ADD_3569 replaced by ADD_4226

//ADD_3568 replaced by ADD_5756

//ADD_3567 replaced by ADD_5756

//ADD_3574 replaced by ADD_4231

//ADD_3573 replaced by ADD_5756

//ADD_3572 replaced by ADD_5756

//ADD_3571 replaced by ADD_5756

//ADD_3570 replaced by ADD_5756

//ADD_3580 replaced by ADD_4237

//ADD_3579 replaced by ADD_5756

//ADD_3578 replaced by ADD_5756

//ADD_3577 replaced by ADD_5756

//ADD_3576 replaced by ADD_5756

//ADD_3575 replaced by ADD_5756

//ADD_3586 replaced by ADD_11592

//ADD_3585 replaced by ADD_5756

//ADD_3584 replaced by ADD_5756

//ADD_3583 replaced by ADD_5756

//ADD_3582 replaced by ADD_5756

//ADD_3581 replaced by ADD_5756

//BADD_1288 replaced by BADD_1312

//BADD_1287 replaced by BADD_1311

//BADD_1286 replaced by BADD_1310

//ADD_3594 replaced by ADD_11602

//ADD_3593 replaced by ADD_11602

//ADD_3592 replaced by ADD_11602

//ADD_3591 replaced by ADD_11602

//ADD_3590 replaced by ADD_11602

//ADD_3589 replaced by ADD_11602

//ADD_3588 replaced by ADD_11602

//ADD_3587 replaced by ADD_11602

//KaratsubaCore_122 replaced by KaratsubaCore_143

//KaratsubaCore_121 replaced by KaratsubaCore_142

//KaratsubaCore_120 replaced by KaratsubaCore_141

//BADD_1291 replaced by BADD_1312

//BADD_1290 replaced by BADD_1311

//BADD_1289 replaced by BADD_1310

//ADD_3602 replaced by ADD_11602

//ADD_3601 replaced by ADD_11602

//ADD_3600 replaced by ADD_11602

//ADD_3599 replaced by ADD_11602

//ADD_3598 replaced by ADD_11602

//ADD_3597 replaced by ADD_11602

//ADD_3596 replaced by ADD_11602

//ADD_3595 replaced by ADD_11602

//KaratsubaCore_125 replaced by KaratsubaCore_143

//KaratsubaCore_124 replaced by KaratsubaCore_142

//KaratsubaCore_123 replaced by KaratsubaCore_141

//BADD_1292 replaced by BADD_1306

//ADD_3608 replaced by ADD_5761

//ADD_3607 replaced by ADD_5756

//ADD_3606 replaced by ADD_5756

//ADD_3605 replaced by ADD_5756

//ADD_3604 replaced by ADD_5756

//ADD_3603 replaced by ADD_5756

//ADD_3614 replaced by ADD_4223

//ADD_3613 replaced by ADD_5756

//ADD_3612 replaced by ADD_5756

//ADD_3611 replaced by ADD_5756

//ADD_3610 replaced by ADD_5756

//ADD_3609 replaced by ADD_5756

//ADD_3616 replaced by ADD_4223

//ADD_3615 replaced by ADD_4226

//ADD_3617 replaced by ADD_4055

//ADD_3618 replaced by ADD_4057

//ADD_3620 replaced by ADD_4223

//ADD_3619 replaced by ADD_4057

//ADD_3621 replaced by ADD_4223

//ADD_3622 replaced by ADD_4060

//ADD_3624 replaced by ADD_4223

//ADD_3623 replaced by ADD_11560

//ADD_3626 replaced by ADD_4223

//ADD_3625 replaced by ADD_4196

//ADD_3628 replaced by ADD_4223

//ADD_3627 replaced by ADD_4132

//ADD_3630 replaced by ADD_4223

//ADD_3629 replaced by ADD_4067

//ADD_3634 replaced by ADD_4223

//ADD_3633 replaced by ADD_5756

//ADD_3632 replaced by ADD_5756

//ADD_3631 replaced by ADD_11592

//ADD_3637 replaced by ADD_4223

//ADD_3636 replaced by ADD_5756

//ADD_3635 replaced by ADD_4168

//ADD_3640 replaced by ADD_4223

//ADD_3639 replaced by ADD_5756

//ADD_3638 replaced by ADD_4076

//ADD_3643 replaced by ADD_4223

//ADD_3642 replaced by ADD_5756

//ADD_3641 replaced by ADD_11592

//ADD_3646 replaced by ADD_4223

//ADD_3645 replaced by ADD_5756

//ADD_3644 replaced by ADD_4106

//ADD_3649 replaced by ADD_4223

//ADD_3648 replaced by ADD_5756

//ADD_3647 replaced by ADD_4085

//ADD_3652 replaced by ADD_4223

//ADD_3651 replaced by ADD_5756

//ADD_3650 replaced by ADD_4158

//ADD_3655 replaced by ADD_4223

//ADD_3654 replaced by ADD_5756

//ADD_3653 replaced by ADD_4091

//ADD_3659 replaced by ADD_4223

//ADD_3658 replaced by ADD_5756

//ADD_3657 replaced by ADD_5756

//ADD_3656 replaced by ADD_4094

//ADD_3663 replaced by ADD_4223

//ADD_3662 replaced by ADD_5756

//ADD_3661 replaced by ADD_5756

//ADD_3660 replaced by ADD_4145

//ADD_3667 replaced by ADD_4223

//ADD_3666 replaced by ADD_5756

//ADD_3665 replaced by ADD_5756

//ADD_3664 replaced by ADD_4212

//ADD_3671 replaced by ADD_4223

//ADD_3670 replaced by ADD_5756

//ADD_3669 replaced by ADD_5756

//ADD_3668 replaced by ADD_4106

//ADD_3676 replaced by ADD_4223

//ADD_3675 replaced by ADD_5756

//ADD_3674 replaced by ADD_5756

//ADD_3673 replaced by ADD_5756

//ADD_3672 replaced by ADD_4212

//ADD_3680 replaced by ADD_4223

//ADD_3679 replaced by ADD_5756

//ADD_3678 replaced by ADD_5756

//ADD_3677 replaced by ADD_4115

//ADD_3685 replaced by ADD_4223

//ADD_3684 replaced by ADD_5756

//ADD_3683 replaced by ADD_5756

//ADD_3682 replaced by ADD_5756

//ADD_3681 replaced by ADD_4231

//ADD_3686 replaced by ADD_11560

//ADD_3689 replaced by ADD_4223

//ADD_3688 replaced by ADD_5756

//ADD_3687 replaced by ADD_4125

//ADD_3691 replaced by ADD_4223

//ADD_3690 replaced by ADD_4131

//ADD_3692 replaced by ADD_4150

//ADD_3693 replaced by ADD_4131

//ADD_3694 replaced by ADD_4132

//ADD_3695 replaced by ADD_4196

//ADD_3696 replaced by ADD_4134

//ADD_3697 replaced by ADD_4139

//ADD_3698 replaced by ADD_4136

//ADD_3700 replaced by ADD_4223

//ADD_3699 replaced by ADD_4172

//ADD_3702 replaced by ADD_4223

//ADD_3701 replaced by ADD_4139

//ADD_3704 replaced by ADD_4223

//ADD_3703 replaced by ADD_4141

//ADD_3706 replaced by ADD_4223

//ADD_3705 replaced by ADD_11602

//ADD_3709 replaced by ADD_4223

//ADD_3708 replaced by ADD_5756

//ADD_3707 replaced by ADD_4145

//ADD_3711 replaced by ADD_4223

//ADD_3710 replaced by ADD_5761

//ADD_3714 replaced by ADD_4223

//ADD_3713 replaced by ADD_5756

//ADD_3712 replaced by ADD_4150

//ADD_3719 replaced by ADD_4223

//ADD_3718 replaced by ADD_5756

//ADD_3717 replaced by ADD_5756

//ADD_3716 replaced by ADD_5756

//ADD_3715 replaced by ADD_4153

//ADD_3723 replaced by ADD_4223

//ADD_3722 replaced by ADD_5756

//ADD_3721 replaced by ADD_5756

//ADD_3720 replaced by ADD_4158

//ADD_3726 replaced by ADD_4223

//ADD_3725 replaced by ADD_5756

//ADD_3724 replaced by ADD_4162

//ADD_3729 replaced by ADD_4223

//ADD_3728 replaced by ADD_5756

//ADD_3727 replaced by ADD_11602

//ADD_3733 replaced by ADD_4223

//ADD_3732 replaced by ADD_5756

//ADD_3731 replaced by ADD_5756

//ADD_3730 replaced by ADD_4168

//ADD_3737 replaced by ADD_4223

//ADD_3736 replaced by ADD_5756

//ADD_3735 replaced by ADD_5756

//ADD_3734 replaced by ADD_4172

//ADD_3741 replaced by ADD_4223

//ADD_3740 replaced by ADD_5756

//ADD_3739 replaced by ADD_5756

//ADD_3738 replaced by ADD_11602

//ADD_3746 replaced by ADD_4223

//ADD_3745 replaced by ADD_5756

//ADD_3744 replaced by ADD_5756

//ADD_3743 replaced by ADD_5756

//ADD_3742 replaced by ADD_11592

//ADD_3752 replaced by ADD_4223

//ADD_3751 replaced by ADD_5756

//ADD_3750 replaced by ADD_5756

//ADD_3749 replaced by ADD_5756

//ADD_3748 replaced by ADD_5756

//ADD_3747 replaced by ADD_11601

//ADD_3757 replaced by ADD_4223

//ADD_3756 replaced by ADD_5756

//ADD_3755 replaced by ADD_5756

//ADD_3754 replaced by ADD_5756

//ADD_3753 replaced by ADD_4191

//ADD_3762 replaced by ADD_4223

//ADD_3761 replaced by ADD_5756

//ADD_3760 replaced by ADD_5756

//ADD_3759 replaced by ADD_5756

//ADD_3758 replaced by ADD_4196

//ADD_3767 replaced by ADD_4223

//ADD_3766 replaced by ADD_5756

//ADD_3765 replaced by ADD_5756

//ADD_3764 replaced by ADD_5756

//ADD_3763 replaced by ADD_4201

//ADD_3773 replaced by ADD_4223

//ADD_3772 replaced by ADD_5756

//ADD_3771 replaced by ADD_5756

//ADD_3770 replaced by ADD_5756

//ADD_3769 replaced by ADD_5756

//ADD_3768 replaced by ADD_4237

//ADD_3779 replaced by ADD_4223

//ADD_3778 replaced by ADD_5756

//ADD_3777 replaced by ADD_5756

//ADD_3776 replaced by ADD_5756

//ADD_3775 replaced by ADD_5756

//ADD_3774 replaced by ADD_4212

//ADD_3785 replaced by ADD_4223

//ADD_3784 replaced by ADD_5756

//ADD_3783 replaced by ADD_5756

//ADD_3782 replaced by ADD_5756

//ADD_3781 replaced by ADD_5756

//ADD_3780 replaced by ADD_4218

//ADD_3788 replaced by ADD_4226

//ADD_3787 replaced by ADD_5756

//ADD_3786 replaced by ADD_5756

//ADD_3793 replaced by ADD_4231

//ADD_3792 replaced by ADD_5756

//ADD_3791 replaced by ADD_5756

//ADD_3790 replaced by ADD_5756

//ADD_3789 replaced by ADD_5756

//ADD_3799 replaced by ADD_4237

//ADD_3798 replaced by ADD_5756

//ADD_3797 replaced by ADD_5756

//ADD_3796 replaced by ADD_5756

//ADD_3795 replaced by ADD_5756

//ADD_3794 replaced by ADD_5756

//ADD_3805 replaced by ADD_11592

//ADD_3804 replaced by ADD_5756

//ADD_3803 replaced by ADD_5756

//ADD_3802 replaced by ADD_5756

//ADD_3801 replaced by ADD_5756

//ADD_3800 replaced by ADD_5756

//BADD_1295 replaced by BADD_1312

//BADD_1294 replaced by BADD_1311

//BADD_1293 replaced by BADD_1310

//ADD_3813 replaced by ADD_11602

//ADD_3812 replaced by ADD_11602

//ADD_3811 replaced by ADD_11602

//ADD_3810 replaced by ADD_11602

//ADD_3809 replaced by ADD_11602

//ADD_3808 replaced by ADD_11602

//ADD_3807 replaced by ADD_11602

//ADD_3806 replaced by ADD_11602

//KaratsubaCore_128 replaced by KaratsubaCore_143

//KaratsubaCore_127 replaced by KaratsubaCore_142

//KaratsubaCore_126 replaced by KaratsubaCore_141

//BADD_1298 replaced by BADD_1312

//BADD_1297 replaced by BADD_1311

//BADD_1296 replaced by BADD_1310

//ADD_3821 replaced by ADD_11602

//ADD_3820 replaced by ADD_11602

//ADD_3819 replaced by ADD_11602

//ADD_3818 replaced by ADD_11602

//ADD_3817 replaced by ADD_11602

//ADD_3816 replaced by ADD_11602

//ADD_3815 replaced by ADD_11602

//ADD_3814 replaced by ADD_11602

//KaratsubaCore_131 replaced by KaratsubaCore_143

//KaratsubaCore_130 replaced by KaratsubaCore_142

//KaratsubaCore_129 replaced by KaratsubaCore_141

//BADD_1299 replaced by BADD_1306

//ADD_3827 replaced by ADD_5761

//ADD_3826 replaced by ADD_5756

//ADD_3825 replaced by ADD_5756

//ADD_3824 replaced by ADD_5756

//ADD_3823 replaced by ADD_5756

//ADD_3822 replaced by ADD_5756

//ADD_3833 replaced by ADD_4223

//ADD_3832 replaced by ADD_5756

//ADD_3831 replaced by ADD_5756

//ADD_3830 replaced by ADD_5756

//ADD_3829 replaced by ADD_5756

//ADD_3828 replaced by ADD_5756

//ADD_3835 replaced by ADD_4223

//ADD_3834 replaced by ADD_4226

//ADD_3836 replaced by ADD_4055

//ADD_3837 replaced by ADD_4057

//ADD_3839 replaced by ADD_4223

//ADD_3838 replaced by ADD_4057

//ADD_3840 replaced by ADD_4223

//ADD_3841 replaced by ADD_4060

//ADD_3843 replaced by ADD_4223

//ADD_3842 replaced by ADD_11560

//ADD_3845 replaced by ADD_4223

//ADD_3844 replaced by ADD_4196

//ADD_3847 replaced by ADD_4223

//ADD_3846 replaced by ADD_4132

//ADD_3849 replaced by ADD_4223

//ADD_3848 replaced by ADD_4067

//ADD_3853 replaced by ADD_4223

//ADD_3852 replaced by ADD_5756

//ADD_3851 replaced by ADD_5756

//ADD_3850 replaced by ADD_11592

//ADD_3856 replaced by ADD_4223

//ADD_3855 replaced by ADD_5756

//ADD_3854 replaced by ADD_4168

//ADD_3859 replaced by ADD_4223

//ADD_3858 replaced by ADD_5756

//ADD_3857 replaced by ADD_4076

//ADD_3862 replaced by ADD_4223

//ADD_3861 replaced by ADD_5756

//ADD_3860 replaced by ADD_11592

//ADD_3865 replaced by ADD_4223

//ADD_3864 replaced by ADD_5756

//ADD_3863 replaced by ADD_4106

//ADD_3868 replaced by ADD_4223

//ADD_3867 replaced by ADD_5756

//ADD_3866 replaced by ADD_4085

//ADD_3871 replaced by ADD_4223

//ADD_3870 replaced by ADD_5756

//ADD_3869 replaced by ADD_4158

//ADD_3874 replaced by ADD_4223

//ADD_3873 replaced by ADD_5756

//ADD_3872 replaced by ADD_4091

//ADD_3878 replaced by ADD_4223

//ADD_3877 replaced by ADD_5756

//ADD_3876 replaced by ADD_5756

//ADD_3875 replaced by ADD_4094

//ADD_3882 replaced by ADD_4223

//ADD_3881 replaced by ADD_5756

//ADD_3880 replaced by ADD_5756

//ADD_3879 replaced by ADD_4145

//ADD_3886 replaced by ADD_4223

//ADD_3885 replaced by ADD_5756

//ADD_3884 replaced by ADD_5756

//ADD_3883 replaced by ADD_4212

//ADD_3890 replaced by ADD_4223

//ADD_3889 replaced by ADD_5756

//ADD_3888 replaced by ADD_5756

//ADD_3887 replaced by ADD_4106

//ADD_3895 replaced by ADD_4223

//ADD_3894 replaced by ADD_5756

//ADD_3893 replaced by ADD_5756

//ADD_3892 replaced by ADD_5756

//ADD_3891 replaced by ADD_4212

//ADD_3899 replaced by ADD_4223

//ADD_3898 replaced by ADD_5756

//ADD_3897 replaced by ADD_5756

//ADD_3896 replaced by ADD_4115

//ADD_3904 replaced by ADD_4223

//ADD_3903 replaced by ADD_5756

//ADD_3902 replaced by ADD_5756

//ADD_3901 replaced by ADD_5756

//ADD_3900 replaced by ADD_4231

//ADD_3905 replaced by ADD_11560

//ADD_3908 replaced by ADD_4223

//ADD_3907 replaced by ADD_5756

//ADD_3906 replaced by ADD_4125

//ADD_3910 replaced by ADD_4223

//ADD_3909 replaced by ADD_4131

//ADD_3911 replaced by ADD_4150

//ADD_3912 replaced by ADD_4131

//ADD_3913 replaced by ADD_4132

//ADD_3914 replaced by ADD_4196

//ADD_3915 replaced by ADD_4134

//ADD_3916 replaced by ADD_4139

//ADD_3917 replaced by ADD_4136

//ADD_3919 replaced by ADD_4223

//ADD_3918 replaced by ADD_4172

//ADD_3921 replaced by ADD_4223

//ADD_3920 replaced by ADD_4139

//ADD_3923 replaced by ADD_4223

//ADD_3922 replaced by ADD_4141

//ADD_3925 replaced by ADD_4223

//ADD_3924 replaced by ADD_11602

//ADD_3928 replaced by ADD_4223

//ADD_3927 replaced by ADD_5756

//ADD_3926 replaced by ADD_4145

//ADD_3930 replaced by ADD_4223

//ADD_3929 replaced by ADD_5761

//ADD_3933 replaced by ADD_4223

//ADD_3932 replaced by ADD_5756

//ADD_3931 replaced by ADD_4150

//ADD_3938 replaced by ADD_4223

//ADD_3937 replaced by ADD_5756

//ADD_3936 replaced by ADD_5756

//ADD_3935 replaced by ADD_5756

//ADD_3934 replaced by ADD_4153

//ADD_3942 replaced by ADD_4223

//ADD_3941 replaced by ADD_5756

//ADD_3940 replaced by ADD_5756

//ADD_3939 replaced by ADD_4158

//ADD_3945 replaced by ADD_4223

//ADD_3944 replaced by ADD_5756

//ADD_3943 replaced by ADD_4162

//ADD_3948 replaced by ADD_4223

//ADD_3947 replaced by ADD_5756

//ADD_3946 replaced by ADD_11602

//ADD_3952 replaced by ADD_4223

//ADD_3951 replaced by ADD_5756

//ADD_3950 replaced by ADD_5756

//ADD_3949 replaced by ADD_4168

//ADD_3956 replaced by ADD_4223

//ADD_3955 replaced by ADD_5756

//ADD_3954 replaced by ADD_5756

//ADD_3953 replaced by ADD_4172

//ADD_3960 replaced by ADD_4223

//ADD_3959 replaced by ADD_5756

//ADD_3958 replaced by ADD_5756

//ADD_3957 replaced by ADD_11602

//ADD_3965 replaced by ADD_4223

//ADD_3964 replaced by ADD_5756

//ADD_3963 replaced by ADD_5756

//ADD_3962 replaced by ADD_5756

//ADD_3961 replaced by ADD_11592

//ADD_3971 replaced by ADD_4223

//ADD_3970 replaced by ADD_5756

//ADD_3969 replaced by ADD_5756

//ADD_3968 replaced by ADD_5756

//ADD_3967 replaced by ADD_5756

//ADD_3966 replaced by ADD_11601

//ADD_3976 replaced by ADD_4223

//ADD_3975 replaced by ADD_5756

//ADD_3974 replaced by ADD_5756

//ADD_3973 replaced by ADD_5756

//ADD_3972 replaced by ADD_4191

//ADD_3981 replaced by ADD_4223

//ADD_3980 replaced by ADD_5756

//ADD_3979 replaced by ADD_5756

//ADD_3978 replaced by ADD_5756

//ADD_3977 replaced by ADD_4196

//ADD_3986 replaced by ADD_4223

//ADD_3985 replaced by ADD_5756

//ADD_3984 replaced by ADD_5756

//ADD_3983 replaced by ADD_5756

//ADD_3982 replaced by ADD_4201

//ADD_3992 replaced by ADD_4223

//ADD_3991 replaced by ADD_5756

//ADD_3990 replaced by ADD_5756

//ADD_3989 replaced by ADD_5756

//ADD_3988 replaced by ADD_5756

//ADD_3987 replaced by ADD_4237

//ADD_3998 replaced by ADD_4223

//ADD_3997 replaced by ADD_5756

//ADD_3996 replaced by ADD_5756

//ADD_3995 replaced by ADD_5756

//ADD_3994 replaced by ADD_5756

//ADD_3993 replaced by ADD_4212

//ADD_4004 replaced by ADD_4223

//ADD_4003 replaced by ADD_5756

//ADD_4002 replaced by ADD_5756

//ADD_4001 replaced by ADD_5756

//ADD_4000 replaced by ADD_5756

//ADD_3999 replaced by ADD_4218

//ADD_4007 replaced by ADD_4226

//ADD_4006 replaced by ADD_5756

//ADD_4005 replaced by ADD_5756

//ADD_4012 replaced by ADD_4231

//ADD_4011 replaced by ADD_5756

//ADD_4010 replaced by ADD_5756

//ADD_4009 replaced by ADD_5756

//ADD_4008 replaced by ADD_5756

//ADD_4018 replaced by ADD_4237

//ADD_4017 replaced by ADD_5756

//ADD_4016 replaced by ADD_5756

//ADD_4015 replaced by ADD_5756

//ADD_4014 replaced by ADD_5756

//ADD_4013 replaced by ADD_5756

//ADD_4024 replaced by ADD_11592

//ADD_4023 replaced by ADD_5756

//ADD_4022 replaced by ADD_5756

//ADD_4021 replaced by ADD_5756

//ADD_4020 replaced by ADD_5756

//ADD_4019 replaced by ADD_5756

//BADD_1302 replaced by BADD_1312

//BADD_1301 replaced by BADD_1311

//BADD_1300 replaced by BADD_1310

//ADD_4032 replaced by ADD_11602

//ADD_4031 replaced by ADD_11602

//ADD_4030 replaced by ADD_11602

//ADD_4029 replaced by ADD_11602

//ADD_4028 replaced by ADD_11602

//ADD_4027 replaced by ADD_11602

//ADD_4026 replaced by ADD_11602

//ADD_4025 replaced by ADD_11602

//KaratsubaCore_134 replaced by KaratsubaCore_143

//KaratsubaCore_133 replaced by KaratsubaCore_142

//KaratsubaCore_132 replaced by KaratsubaCore_141

//BADD_1305 replaced by BADD_1312

//BADD_1304 replaced by BADD_1311

//BADD_1303 replaced by BADD_1310

//ADD_4040 replaced by ADD_11602

//ADD_4039 replaced by ADD_11602

//ADD_4038 replaced by ADD_11602

//ADD_4037 replaced by ADD_11602

//ADD_4036 replaced by ADD_11602

//ADD_4035 replaced by ADD_11602

//ADD_4034 replaced by ADD_11602

//ADD_4033 replaced by ADD_11602

//KaratsubaCore_137 replaced by KaratsubaCore_143

//KaratsubaCore_136 replaced by KaratsubaCore_142

//KaratsubaCore_135 replaced by KaratsubaCore_141

module BADD_1306 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  input               io_c,
  output     [378:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [63:0]   adder_adds_0_io_A_0;
  wire       [63:0]   adder_adds_0_io_A_1;
  wire       [63:0]   adder_adds_1_io_A_0;
  wire       [63:0]   adder_adds_1_io_A_1;
  wire       [63:0]   adder_adds_2_io_A_0;
  wire       [63:0]   adder_adds_2_io_A_1;
  wire       [63:0]   adder_adds_3_io_A_0;
  wire       [63:0]   adder_adds_3_io_A_1;
  wire       [63:0]   adder_adds_4_io_A_0;
  wire       [63:0]   adder_adds_4_io_A_1;
  wire       [57:0]   adder_adds_5_io_A_0;
  wire       [57:0]   adder_adds_5_io_A_1;
  wire       [64:0]   adder_adds_0_io_S;
  wire       [64:0]   adder_adds_1_io_S;
  wire       [64:0]   adder_adds_2_io_S;
  wire       [64:0]   adder_adds_3_io_S;
  wire       [64:0]   adder_adds_4_io_S;
  wire       [58:0]   adder_adds_5_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  reg        [57:0]   _zz_io_s_21;

  ADD_5756 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[63:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[64:0]  )  //o
  );
  ADD_5756 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[63:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[63:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[64:0]  )  //o
  );
  ADD_5761 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[57:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[57:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[58:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[63 : 0];
  assign adder_adds_1_io_A_0 = io_a[127 : 64];
  assign adder_adds_2_io_A_0 = io_a[191 : 128];
  assign adder_adds_3_io_A_0 = io_a[255 : 192];
  assign adder_adds_4_io_A_0 = io_a[319 : 256];
  assign adder_adds_5_io_A_0 = io_a[377 : 320];
  assign adder_adds_0_io_A_1 = io_b[63 : 0];
  assign adder_adds_1_io_A_1 = io_b[127 : 64];
  assign adder_adds_2_io_A_1 = io_b[191 : 128];
  assign adder_adds_3_io_A_1 = io_b[255 : 192];
  assign adder_adds_4_io_A_1 = io_b[319 : 256];
  assign adder_adds_5_io_A_1 = io_b[377 : 320];
  assign io_s = {_zz_io_s,{_zz_io_s_21,{_zz_io_s_20,{_zz_io_s_18,{_zz_io_s_15,{_zz_io_s_11,_zz_io_s_6}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[64];
    _zz_io_CIN_1 <= adder_adds_1_io_S[64];
    _zz_io_CIN_2 <= adder_adds_2_io_S[64];
    _zz_io_CIN_3 <= adder_adds_3_io_S[64];
    _zz_io_CIN_4 <= adder_adds_4_io_S[64];
    _zz_io_s <= adder_adds_5_io_S[58];
    _zz_io_s_1 <= adder_adds_0_io_S[63 : 0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= adder_adds_1_io_S[63 : 0];
    _zz_io_s_8 <= _zz_io_s_7;
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= adder_adds_2_io_S[63 : 0];
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= adder_adds_3_io_S[63 : 0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= adder_adds_4_io_S[63 : 0];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_21 <= adder_adds_5_io_S[57 : 0];
  end


endmodule

//ADD_4046 replaced by ADD_5761

//ADD_4045 replaced by ADD_5756

//ADD_4044 replaced by ADD_5756

//ADD_4043 replaced by ADD_5756

//ADD_4042 replaced by ADD_5756

//ADD_4041 replaced by ADD_5756

//ADD_4052 replaced by ADD_4223

//ADD_4051 replaced by ADD_5756

//ADD_4050 replaced by ADD_5756

//ADD_4049 replaced by ADD_5756

//ADD_4048 replaced by ADD_5756

//ADD_4047 replaced by ADD_5756

//ADD_4054 replaced by ADD_4223

//ADD_4053 replaced by ADD_4226

module ADD_4055 (
  input      [36:0]   io_A_0,
  input      [36:0]   io_A_1,
  input               io_CIN,
  output     [37:0]   io_S
);

  wire       [37:0]   _zz_io_S;
  wire       [37:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {37'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4056 replaced by ADD_4057

//ADD_4058 replaced by ADD_4223

module ADD_4057 (
  input      [9:0]    io_A_0,
  input      [9:0]    io_A_1,
  input               io_CIN,
  output     [10:0]   io_S
);

  wire       [10:0]   _zz_io_S;
  wire       [10:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {10'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4059 replaced by ADD_4223

module ADD_4060 (
  input      [54:0]   io_A_0,
  input      [54:0]   io_A_1,
  input               io_CIN,
  output     [55:0]   io_S
);

  wire       [55:0]   _zz_io_S;
  wire       [55:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {55'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4062 replaced by ADD_4223

//ADD_4061 replaced by ADD_11560

//ADD_4064 replaced by ADD_4223

//ADD_4063 replaced by ADD_4196

//ADD_4066 replaced by ADD_4223

//ADD_4065 replaced by ADD_4132

//ADD_4068 replaced by ADD_4223

module ADD_4067 (
  input      [37:0]   io_A_0,
  input      [37:0]   io_A_1,
  input               io_CIN,
  output     [38:0]   io_S
);

  wire       [38:0]   _zz_io_S;
  wire       [38:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {38'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4072 replaced by ADD_4223

//ADD_4071 replaced by ADD_5756

//ADD_4070 replaced by ADD_5756

//ADD_4069 replaced by ADD_11592

//ADD_4075 replaced by ADD_4223

//ADD_4074 replaced by ADD_5756

//ADD_4073 replaced by ADD_4168

//ADD_4078 replaced by ADD_4223

//ADD_4077 replaced by ADD_5756

module ADD_4076 (
  input      [6:0]    io_A_0,
  input      [6:0]    io_A_1,
  input               io_CIN,
  output     [7:0]    io_S
);

  wire       [7:0]    _zz_io_S;
  wire       [7:0]    _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {7'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4081 replaced by ADD_4223

//ADD_4080 replaced by ADD_5756

//ADD_4079 replaced by ADD_11592

//ADD_4084 replaced by ADD_4223

//ADD_4083 replaced by ADD_5756

//ADD_4082 replaced by ADD_4106

//ADD_4087 replaced by ADD_4223

//ADD_4086 replaced by ADD_5756

module ADD_4085 (
  input      [43:0]   io_A_0,
  input      [43:0]   io_A_1,
  input               io_CIN,
  output     [44:0]   io_S
);

  wire       [44:0]   _zz_io_S;
  wire       [44:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {44'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4090 replaced by ADD_4223

//ADD_4089 replaced by ADD_5756

//ADD_4088 replaced by ADD_4158

//ADD_4093 replaced by ADD_4223

//ADD_4092 replaced by ADD_5756

module ADD_4091 (
  input      [59:0]   io_A_0,
  input      [59:0]   io_A_1,
  input               io_CIN,
  output     [60:0]   io_S
);

  wire       [60:0]   _zz_io_S;
  wire       [60:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {60'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4097 replaced by ADD_4223

//ADD_4096 replaced by ADD_5756

//ADD_4095 replaced by ADD_5756

module ADD_4094 (
  input      [33:0]   io_A_0,
  input      [33:0]   io_A_1,
  input               io_CIN,
  output     [34:0]   io_S
);

  wire       [34:0]   _zz_io_S;
  wire       [34:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {34'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4101 replaced by ADD_4223

//ADD_4100 replaced by ADD_5756

//ADD_4099 replaced by ADD_5756

//ADD_4098 replaced by ADD_4145

//ADD_4105 replaced by ADD_4223

//ADD_4104 replaced by ADD_5756

//ADD_4103 replaced by ADD_5756

//ADD_4102 replaced by ADD_4212

//ADD_4109 replaced by ADD_4223

//ADD_4108 replaced by ADD_5756

//ADD_4107 replaced by ADD_5756

module ADD_4106 (
  input      [18:0]   io_A_0,
  input      [18:0]   io_A_1,
  input               io_CIN,
  output     [19:0]   io_S
);

  wire       [19:0]   _zz_io_S;
  wire       [19:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {19'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4114 replaced by ADD_4223

//ADD_4113 replaced by ADD_5756

//ADD_4112 replaced by ADD_5756

//ADD_4111 replaced by ADD_5756

//ADD_4110 replaced by ADD_4212

//ADD_4118 replaced by ADD_4223

//ADD_4117 replaced by ADD_5756

//ADD_4116 replaced by ADD_5756

module ADD_4115 (
  input      [38:0]   io_A_0,
  input      [38:0]   io_A_1,
  input               io_CIN,
  output     [39:0]   io_S
);

  wire       [39:0]   _zz_io_S;
  wire       [39:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {39'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4123 replaced by ADD_4223

//ADD_4122 replaced by ADD_5756

//ADD_4121 replaced by ADD_5756

//ADD_4120 replaced by ADD_5756

//ADD_4119 replaced by ADD_4231

//ADD_4124 replaced by ADD_11560

//ADD_4127 replaced by ADD_4223

//ADD_4126 replaced by ADD_5756

module ADD_4125 (
  input      [39:0]   io_A_0,
  input      [39:0]   io_A_1,
  input               io_CIN,
  output     [40:0]   io_S
);

  wire       [40:0]   _zz_io_S;
  wire       [40:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {40'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4129 replaced by ADD_4223

//ADD_4128 replaced by ADD_4131

//ADD_4130 replaced by ADD_4150

module ADD_4131 (
  input      [20:0]   io_A_0,
  input      [20:0]   io_A_1,
  input               io_CIN,
  output     [21:0]   io_S
);

  wire       [21:0]   _zz_io_S;
  wire       [21:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {21'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

module ADD_4132 (
  input      [15:0]   io_A_0,
  input      [15:0]   io_A_1,
  input               io_CIN,
  output     [16:0]   io_S
);

  wire       [16:0]   _zz_io_S;
  wire       [16:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {16'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4133 replaced by ADD_4196

module ADD_4134 (
  input      [46:0]   io_A_0,
  input      [46:0]   io_A_1,
  input               io_CIN,
  output     [47:0]   io_S
);

  wire       [47:0]   _zz_io_S;
  wire       [47:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {47'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4135 replaced by ADD_4139

module ADD_4136 (
  input      [50:0]   io_A_0,
  input      [50:0]   io_A_1,
  input               io_CIN,
  output     [51:0]   io_S
);

  wire       [51:0]   _zz_io_S;
  wire       [51:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {51'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4138 replaced by ADD_4223

//ADD_4137 replaced by ADD_4172

//ADD_4140 replaced by ADD_4223

module ADD_4139 (
  input      [42:0]   io_A_0,
  input      [42:0]   io_A_1,
  input               io_CIN,
  output     [43:0]   io_S
);

  wire       [43:0]   _zz_io_S;
  wire       [43:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {43'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4142 replaced by ADD_4223

module ADD_4141 (
  input      [32:0]   io_A_0,
  input      [32:0]   io_A_1,
  input               io_CIN,
  output     [33:0]   io_S
);

  wire       [33:0]   _zz_io_S;
  wire       [33:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {33'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4144 replaced by ADD_4223

//ADD_4143 replaced by ADD_11602

//ADD_4147 replaced by ADD_4223

//ADD_4146 replaced by ADD_5756

module ADD_4145 (
  input      [13:0]   io_A_0,
  input      [13:0]   io_A_1,
  input               io_CIN,
  output     [14:0]   io_S
);

  wire       [14:0]   _zz_io_S;
  wire       [14:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {14'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4149 replaced by ADD_4223

//ADD_4148 replaced by ADD_5761

//ADD_4152 replaced by ADD_4223

//ADD_4151 replaced by ADD_5756

module ADD_4150 (
  input      [31:0]   io_A_0,
  input      [31:0]   io_A_1,
  input               io_CIN,
  output     [32:0]   io_S
);

  wire       [32:0]   _zz_io_S;
  wire       [32:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {32'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4157 replaced by ADD_4223

//ADD_4156 replaced by ADD_5756

//ADD_4155 replaced by ADD_5756

//ADD_4154 replaced by ADD_5756

module ADD_4153 (
  input      [11:0]   io_A_0,
  input      [11:0]   io_A_1,
  input               io_CIN,
  output     [12:0]   io_S
);

  wire       [12:0]   _zz_io_S;
  wire       [12:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {12'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4161 replaced by ADD_4223

//ADD_4160 replaced by ADD_5756

//ADD_4159 replaced by ADD_5756

module ADD_4158 (
  input      [27:0]   io_A_0,
  input      [27:0]   io_A_1,
  input               io_CIN,
  output     [28:0]   io_S
);

  wire       [28:0]   _zz_io_S;
  wire       [28:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {28'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4164 replaced by ADD_4223

//ADD_4163 replaced by ADD_5756

module ADD_4162 (
  input      [53:0]   io_A_0,
  input      [53:0]   io_A_1,
  input               io_CIN,
  output     [54:0]   io_S
);

  wire       [54:0]   _zz_io_S;
  wire       [54:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {54'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4167 replaced by ADD_4223

//ADD_4166 replaced by ADD_5756

//ADD_4165 replaced by ADD_11602

//ADD_4171 replaced by ADD_4223

//ADD_4170 replaced by ADD_5756

//ADD_4169 replaced by ADD_5756

module ADD_4168 (
  input      [22:0]   io_A_0,
  input      [22:0]   io_A_1,
  input               io_CIN,
  output     [23:0]   io_S
);

  wire       [23:0]   _zz_io_S;
  wire       [23:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {23'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4175 replaced by ADD_4223

//ADD_4174 replaced by ADD_5756

//ADD_4173 replaced by ADD_5756

module ADD_4172 (
  input      [52:0]   io_A_0,
  input      [52:0]   io_A_1,
  input               io_CIN,
  output     [53:0]   io_S
);

  wire       [53:0]   _zz_io_S;
  wire       [53:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {53'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4179 replaced by ADD_4223

//ADD_4178 replaced by ADD_5756

//ADD_4177 replaced by ADD_5756

//ADD_4176 replaced by ADD_11602

//ADD_4184 replaced by ADD_4223

//ADD_4183 replaced by ADD_5756

//ADD_4182 replaced by ADD_5756

//ADD_4181 replaced by ADD_5756

//ADD_4180 replaced by ADD_11592

//ADD_4190 replaced by ADD_4223

//ADD_4189 replaced by ADD_5756

//ADD_4188 replaced by ADD_5756

//ADD_4187 replaced by ADD_5756

//ADD_4186 replaced by ADD_5756

//ADD_4185 replaced by ADD_11601

//ADD_4195 replaced by ADD_4223

//ADD_4194 replaced by ADD_5756

//ADD_4193 replaced by ADD_5756

//ADD_4192 replaced by ADD_5756

module ADD_4191 (
  input      [29:0]   io_A_0,
  input      [29:0]   io_A_1,
  input               io_CIN,
  output     [30:0]   io_S
);

  wire       [30:0]   _zz_io_S;
  wire       [30:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {30'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4200 replaced by ADD_4223

//ADD_4199 replaced by ADD_5756

//ADD_4198 replaced by ADD_5756

//ADD_4197 replaced by ADD_5756

module ADD_4196 (
  input      [25:0]   io_A_0,
  input      [25:0]   io_A_1,
  input               io_CIN,
  output     [26:0]   io_S
);

  wire       [26:0]   _zz_io_S;
  wire       [26:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {26'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4205 replaced by ADD_4223

//ADD_4204 replaced by ADD_5756

//ADD_4203 replaced by ADD_5756

//ADD_4202 replaced by ADD_5756

module ADD_4201 (
  input      [35:0]   io_A_0,
  input      [35:0]   io_A_1,
  input               io_CIN,
  output     [36:0]   io_S
);

  wire       [36:0]   _zz_io_S;
  wire       [36:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {36'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4211 replaced by ADD_4223

//ADD_4210 replaced by ADD_5756

//ADD_4209 replaced by ADD_5756

//ADD_4208 replaced by ADD_5756

//ADD_4207 replaced by ADD_5756

//ADD_4206 replaced by ADD_4237

//ADD_4217 replaced by ADD_4223

//ADD_4216 replaced by ADD_5756

//ADD_4215 replaced by ADD_5756

//ADD_4214 replaced by ADD_5756

//ADD_4213 replaced by ADD_5756

module ADD_4212 (
  input      [7:0]    io_A_0,
  input      [7:0]    io_A_1,
  input               io_CIN,
  output     [8:0]    io_S
);

  wire       [8:0]    _zz_io_S;
  wire       [8:0]    _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {8'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

module ADD_4223 (
  input      [58:0]   io_A_0,
  input      [58:0]   io_A_1,
  input               io_CIN,
  output     [59:0]   io_S
);

  wire       [59:0]   _zz_io_S;
  wire       [59:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {59'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4222 replaced by ADD_5756

//ADD_4221 replaced by ADD_5756

//ADD_4220 replaced by ADD_5756

//ADD_4219 replaced by ADD_5756

module ADD_4218 (
  input      [17:0]   io_A_0,
  input      [17:0]   io_A_1,
  input               io_CIN,
  output     [18:0]   io_S
);

  wire       [18:0]   _zz_io_S;
  wire       [18:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {18'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

module ADD_4226 (
  input      [61:0]   io_A_0,
  input      [61:0]   io_A_1,
  input               io_CIN,
  output     [62:0]   io_S
);

  wire       [62:0]   _zz_io_S;
  wire       [62:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {62'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4225 replaced by ADD_5756

//ADD_4224 replaced by ADD_5756

module ADD_4231 (
  input      [16:0]   io_A_0,
  input      [16:0]   io_A_1,
  input               io_CIN,
  output     [17:0]   io_S
);

  wire       [17:0]   _zz_io_S;
  wire       [17:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {17'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4230 replaced by ADD_5756

//ADD_4229 replaced by ADD_5756

//ADD_4228 replaced by ADD_5756

//ADD_4227 replaced by ADD_5756

module ADD_4237 (
  input      [12:0]   io_A_0,
  input      [12:0]   io_A_1,
  input               io_CIN,
  output     [13:0]   io_S
);

  wire       [13:0]   _zz_io_S;
  wire       [13:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {13'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_4236 replaced by ADD_5756

//ADD_4235 replaced by ADD_5756

//ADD_4234 replaced by ADD_5756

//ADD_4233 replaced by ADD_5756

//ADD_4232 replaced by ADD_5756

//ADD_4243 replaced by ADD_11592

//ADD_4242 replaced by ADD_5756

//ADD_4241 replaced by ADD_5756

//ADD_4240 replaced by ADD_5756

//ADD_4239 replaced by ADD_5756

//ADD_4238 replaced by ADD_5756

//BADD_1309 replaced by BADD_1312

//BADD_1308 replaced by BADD_1311

//BADD_1307 replaced by BADD_1310

//ADD_4251 replaced by ADD_11602

//ADD_4250 replaced by ADD_11602

//ADD_4249 replaced by ADD_11602

//ADD_4248 replaced by ADD_11602

//ADD_4247 replaced by ADD_11602

//ADD_4246 replaced by ADD_11602

//ADD_4245 replaced by ADD_11602

//ADD_4244 replaced by ADD_11602

//KaratsubaCore_140 replaced by KaratsubaCore_143

//KaratsubaCore_139 replaced by KaratsubaCore_142

//KaratsubaCore_138 replaced by KaratsubaCore_141

module BADD_1312 (
  input      [575:0]  io_a,
  input      [575:0]  io_b,
  input               io_c,
  output     [576:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [47:0]   adder_adds_4_io_A_0;
  wire       [47:0]   adder_adds_4_io_A_1;
  wire       [47:0]   adder_adds_5_io_A_0;
  wire       [47:0]   adder_adds_5_io_A_1;
  wire       [47:0]   adder_adds_6_io_A_0;
  wire       [47:0]   adder_adds_6_io_A_1;
  wire       [47:0]   adder_adds_7_io_A_0;
  wire       [47:0]   adder_adds_7_io_A_1;
  wire       [47:0]   adder_adds_8_io_A_0;
  wire       [47:0]   adder_adds_8_io_A_1;
  wire       [47:0]   adder_adds_9_io_A_0;
  wire       [47:0]   adder_adds_9_io_A_1;
  wire       [47:0]   adder_adds_10_io_A_0;
  wire       [47:0]   adder_adds_10_io_A_1;
  wire       [47:0]   adder_adds_11_io_A_0;
  wire       [47:0]   adder_adds_11_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  wire       [48:0]   adder_adds_4_io_S;
  wire       [48:0]   adder_adds_5_io_S;
  wire       [48:0]   adder_adds_6_io_S;
  wire       [48:0]   adder_adds_7_io_S;
  wire       [48:0]   adder_adds_8_io_S;
  wire       [48:0]   adder_adds_9_io_S;
  wire       [48:0]   adder_adds_10_io_S;
  wire       [48:0]   adder_adds_11_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_CIN_5;
  reg                 _zz_io_CIN_6;
  reg                 _zz_io_CIN_7;
  reg                 _zz_io_CIN_8;
  reg                 _zz_io_CIN_9;
  reg                 _zz_io_CIN_10;
  reg                 _zz_io_s;
  reg                 _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [47:0]   _zz_io_s_5;
  reg        [47:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg        [47:0]   _zz_io_s_8;
  reg        [47:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg        [47:0]   _zz_io_s_11;
  reg        [47:0]   _zz_io_s_12;
  reg        [47:0]   _zz_io_s_13;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_6 (
    .io_A_0 (adder_adds_6_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_6_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_5             ), //i
    .io_S   (adder_adds_6_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_7 (
    .io_A_0 (adder_adds_7_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_7_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_6             ), //i
    .io_S   (adder_adds_7_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_8 (
    .io_A_0 (adder_adds_8_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_8_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_7             ), //i
    .io_S   (adder_adds_8_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_9 (
    .io_A_0 (adder_adds_9_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_9_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_8             ), //i
    .io_S   (adder_adds_9_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_10 (
    .io_A_0 (adder_adds_10_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_10_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_9              ), //i
    .io_S   (adder_adds_10_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_11 (
    .io_A_0 (adder_adds_11_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_11_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_10             ), //i
    .io_S   (adder_adds_11_io_S[48:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_4_io_A_0 = io_a[239 : 192];
  assign adder_adds_5_io_A_0 = io_a[287 : 240];
  assign adder_adds_6_io_A_0 = io_a[335 : 288];
  assign adder_adds_7_io_A_0 = io_a[383 : 336];
  assign adder_adds_8_io_A_0 = io_a[431 : 384];
  assign adder_adds_9_io_A_0 = io_a[479 : 432];
  assign adder_adds_10_io_A_0 = io_a[527 : 480];
  assign adder_adds_11_io_A_0 = io_a[575 : 528];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[143 : 96];
  assign adder_adds_3_io_A_1 = io_b[191 : 144];
  assign adder_adds_4_io_A_1 = io_b[239 : 192];
  assign adder_adds_5_io_A_1 = io_b[287 : 240];
  assign adder_adds_6_io_A_1 = io_b[335 : 288];
  assign adder_adds_7_io_A_1 = io_b[383 : 336];
  assign adder_adds_8_io_A_1 = io_b[431 : 384];
  assign adder_adds_9_io_A_1 = io_b[479 : 432];
  assign adder_adds_10_io_A_1 = io_b[527 : 480];
  assign adder_adds_11_io_A_1 = io_b[575 : 528];
  assign io_s = {_zz_io_s_1,{_zz_io_s_13,{_zz_io_s_12,{_zz_io_s_11,{_zz_io_s_10,{_zz_io_s_9,{_zz_io_s_8,{_zz_io_s_7,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,_zz_io_s_2}}}}}}}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_CIN_3 <= adder_adds_3_io_S[48];
    _zz_io_CIN_4 <= adder_adds_4_io_S[48];
    _zz_io_CIN_5 <= adder_adds_5_io_S[48];
    _zz_io_CIN_6 <= adder_adds_6_io_S[48];
    _zz_io_CIN_7 <= adder_adds_7_io_S[48];
    _zz_io_CIN_8 <= adder_adds_8_io_S[48];
    _zz_io_CIN_9 <= adder_adds_9_io_S[48];
    _zz_io_CIN_10 <= adder_adds_10_io_S[48];
    _zz_io_s <= adder_adds_11_io_S[48];
    _zz_io_s_1 <= _zz_io_s;
    _zz_io_s_2 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_3_io_S[47 : 0];
    _zz_io_s_6 <= adder_adds_4_io_S[47 : 0];
    _zz_io_s_7 <= adder_adds_5_io_S[47 : 0];
    _zz_io_s_8 <= adder_adds_6_io_S[47 : 0];
    _zz_io_s_9 <= adder_adds_7_io_S[47 : 0];
    _zz_io_s_10 <= adder_adds_8_io_S[47 : 0];
    _zz_io_s_11 <= adder_adds_9_io_S[47 : 0];
    _zz_io_s_12 <= adder_adds_10_io_S[47 : 0];
    _zz_io_s_13 <= adder_adds_11_io_S[47 : 0];
  end


endmodule

module BADD_1311 (
  input      [384:0]  io_a,
  input      [384:0]  io_b,
  input               io_c,
  output     [385:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [47:0]   adder_adds_4_io_A_0;
  wire       [47:0]   adder_adds_4_io_A_1;
  wire       [47:0]   adder_adds_5_io_A_0;
  wire       [47:0]   adder_adds_5_io_A_1;
  wire       [47:0]   adder_adds_6_io_A_0;
  wire       [47:0]   adder_adds_6_io_A_1;
  wire       [47:0]   adder_adds_7_io_A_0;
  wire       [47:0]   adder_adds_7_io_A_1;
  wire       [0:0]    adder_adds_8_io_A_0;
  wire       [0:0]    adder_adds_8_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  wire       [48:0]   adder_adds_4_io_S;
  wire       [48:0]   adder_adds_5_io_S;
  wire       [48:0]   adder_adds_6_io_S;
  wire       [48:0]   adder_adds_7_io_S;
  wire       [1:0]    adder_adds_8_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_CIN_5;
  reg                 _zz_io_CIN_6;
  reg                 _zz_io_CIN_7;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [47:0]   _zz_io_s_5;
  reg        [47:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg        [47:0]   _zz_io_s_8;
  reg        [0:0]    _zz_io_s_9;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_6 (
    .io_A_0 (adder_adds_6_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_6_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_5             ), //i
    .io_S   (adder_adds_6_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_7 (
    .io_A_0 (adder_adds_7_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_7_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_6             ), //i
    .io_S   (adder_adds_7_io_S[48:0]  )  //o
  );
  ADD_11601 adder_adds_8 (
    .io_A_0 (adder_adds_8_io_A_0   ), //i
    .io_A_1 (adder_adds_8_io_A_1   ), //i
    .io_CIN (_zz_io_CIN_7          ), //i
    .io_S   (adder_adds_8_io_S[1:0])  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_4_io_A_0 = io_a[239 : 192];
  assign adder_adds_5_io_A_0 = io_a[287 : 240];
  assign adder_adds_6_io_A_0 = io_a[335 : 288];
  assign adder_adds_7_io_A_0 = io_a[383 : 336];
  assign adder_adds_8_io_A_0 = io_a[384 : 384];
  assign adder_adds_0_io_A_1 = (~ io_b[47 : 0]);
  assign adder_adds_1_io_A_1 = (~ io_b[95 : 48]);
  assign adder_adds_2_io_A_1 = (~ io_b[143 : 96]);
  assign adder_adds_3_io_A_1 = (~ io_b[191 : 144]);
  assign adder_adds_4_io_A_1 = (~ io_b[239 : 192]);
  assign adder_adds_5_io_A_1 = (~ io_b[287 : 240]);
  assign adder_adds_6_io_A_1 = (~ io_b[335 : 288]);
  assign adder_adds_7_io_A_1 = (~ io_b[383 : 336]);
  assign adder_adds_8_io_A_1 = (~ io_b[384 : 384]);
  assign io_s = {_zz_io_s,{_zz_io_s_9,{_zz_io_s_8,{_zz_io_s_7,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_CIN_3 <= adder_adds_3_io_S[48];
    _zz_io_CIN_4 <= adder_adds_4_io_S[48];
    _zz_io_CIN_5 <= adder_adds_5_io_S[48];
    _zz_io_CIN_6 <= adder_adds_6_io_S[48];
    _zz_io_CIN_7 <= adder_adds_7_io_S[48];
    _zz_io_s <= (! adder_adds_8_io_S[1]);
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[47 : 0];
    _zz_io_s_6 <= adder_adds_5_io_S[47 : 0];
    _zz_io_s_7 <= adder_adds_6_io_S[47 : 0];
    _zz_io_s_8 <= adder_adds_7_io_S[47 : 0];
    _zz_io_s_9 <= adder_adds_8_io_S[0 : 0];
  end


endmodule

module BADD_1310 (
  input      [383:0]  io_a,
  input      [383:0]  io_b,
  input               io_c,
  output     [384:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [47:0]   adder_adds_4_io_A_0;
  wire       [47:0]   adder_adds_4_io_A_1;
  wire       [47:0]   adder_adds_5_io_A_0;
  wire       [47:0]   adder_adds_5_io_A_1;
  wire       [47:0]   adder_adds_6_io_A_0;
  wire       [47:0]   adder_adds_6_io_A_1;
  wire       [47:0]   adder_adds_7_io_A_0;
  wire       [47:0]   adder_adds_7_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  wire       [48:0]   adder_adds_4_io_S;
  wire       [48:0]   adder_adds_5_io_S;
  wire       [48:0]   adder_adds_6_io_S;
  wire       [48:0]   adder_adds_7_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_CIN_5;
  reg                 _zz_io_CIN_6;
  reg                 _zz_io_s;
  reg                 _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [47:0]   _zz_io_s_5;
  reg        [47:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg        [47:0]   _zz_io_s_8;
  reg        [47:0]   _zz_io_s_9;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_6 (
    .io_A_0 (adder_adds_6_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_6_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_5             ), //i
    .io_S   (adder_adds_6_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_7 (
    .io_A_0 (adder_adds_7_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_7_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_6             ), //i
    .io_S   (adder_adds_7_io_S[48:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_4_io_A_0 = io_a[239 : 192];
  assign adder_adds_5_io_A_0 = io_a[287 : 240];
  assign adder_adds_6_io_A_0 = io_a[335 : 288];
  assign adder_adds_7_io_A_0 = io_a[383 : 336];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[143 : 96];
  assign adder_adds_3_io_A_1 = io_b[191 : 144];
  assign adder_adds_4_io_A_1 = io_b[239 : 192];
  assign adder_adds_5_io_A_1 = io_b[287 : 240];
  assign adder_adds_6_io_A_1 = io_b[335 : 288];
  assign adder_adds_7_io_A_1 = io_b[383 : 336];
  assign io_s = {_zz_io_s_1,{_zz_io_s_9,{_zz_io_s_8,{_zz_io_s_7,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,_zz_io_s_2}}}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_CIN_3 <= adder_adds_3_io_S[48];
    _zz_io_CIN_4 <= adder_adds_4_io_S[48];
    _zz_io_CIN_5 <= adder_adds_5_io_S[48];
    _zz_io_CIN_6 <= adder_adds_6_io_S[48];
    _zz_io_s <= adder_adds_7_io_S[48];
    _zz_io_s_1 <= _zz_io_s;
    _zz_io_s_2 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_3_io_S[47 : 0];
    _zz_io_s_6 <= adder_adds_4_io_S[47 : 0];
    _zz_io_s_7 <= adder_adds_5_io_S[47 : 0];
    _zz_io_s_8 <= adder_adds_6_io_S[47 : 0];
    _zz_io_s_9 <= adder_adds_7_io_S[47 : 0];
  end


endmodule

//ADD_4259 replaced by ADD_11602

//ADD_4258 replaced by ADD_11602

//ADD_4257 replaced by ADD_11602

//ADD_4256 replaced by ADD_11602

//ADD_4255 replaced by ADD_11602

//ADD_4254 replaced by ADD_11602

//ADD_4253 replaced by ADD_11602

//ADD_4252 replaced by ADD_11602

module KaratsubaCore_143 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_a_2,
  input      [47:0]   io_a_3,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  input      [47:0]   io_b_2,
  input      [47:0]   io_b_3,
  output reg [383:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [192:0]  karatsuba_add2_io_a;
  wire       [287:0]  karatsuba_noExtend_add3_io_a;
  reg        [287:0]  karatsuba_noExtend_add3_io_b;
  wire       [191:0]  karatsuba_lsbMul_io_p;
  wire       [193:0]  karatsuba_midMul_io_p;
  wire       [191:0]  karatsuba_msbMul_io_p;
  wire       [48:0]   karatsuba_midAdd_0_0_io_S;
  wire       [48:0]   karatsuba_midAdd_0_1_io_S;
  wire       [48:0]   karatsuba_midAdd_1_0_io_S;
  wire       [48:0]   karatsuba_midAdd_1_1_io_S;
  wire       [192:0]  karatsuba_add1_io_s;
  wire       [193:0]  karatsuba_add2_io_s;
  wire       [288:0]  karatsuba_noExtend_add3_io_s;
  wire       [192:0]  _zz_io_a;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_a_1;
  reg        [48:0]   _zz_io_b_0;
  reg        [48:0]   _zz_io_b_1;
  reg        [192:0]  karatsuba_msbMul_karatsuba_add1_io_s_delay_1;
  reg        [95:0]   _zz_io_b;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_5;
  reg        [95:0]   _zz_io_p;
  reg        [95:0]   _zz_io_p_1;

  assign _zz_io_a = karatsuba_add2_io_s[192:0];
  KaratsubaCore_465 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]                ), //i
    .io_a_1 (io_a_1[47:0]                ), //i
    .io_b_0 (io_b_0[47:0]                ), //i
    .io_b_1 (io_b_1[47:0]                ), //i
    .io_p   (karatsuba_lsbMul_io_p[191:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_466 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]            ), //i
    .io_a_1 (_zz_io_a_1[48:0]            ), //i
    .io_b_0 (_zz_io_b_0[48:0]            ), //i
    .io_b_1 (_zz_io_b_1[48:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[193:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_467 karatsuba_msbMul (
    .io_a_0 (io_a_2[47:0]                ), //i
    .io_a_1 (io_a_3[47:0]                ), //i
    .io_b_0 (io_b_2[47:0]                ), //i
    .io_b_1 (io_b_3[47:0]                ), //i
    .io_p   (karatsuba_msbMul_io_p[191:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  ADD_11602 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[47:0]                   ), //i
    .io_A_1 (io_a_2[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_0_1 (
    .io_A_0 (io_a_1[47:0]                   ), //i
    .io_A_1 (io_a_3[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_1_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[47:0]                   ), //i
    .io_A_1 (io_b_2[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_1 (
    .io_A_0 (io_b_1[47:0]                   ), //i
    .io_A_1 (io_b_3[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_1_io_S[48:0])  //o
  );
  BADD_1670 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[191:0]), //i
    .io_b   (karatsuba_msbMul_io_p[191:0]), //i
    .io_c   (1'b0                        ), //i
    .io_s   (karatsuba_add1_io_s[192:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_1671 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[192:0]                         ), //i
    .io_b   (karatsuba_msbMul_karatsuba_add1_io_s_delay_1[192:0]), //i
    .io_c   (1'b1                                               ), //i
    .io_s   (karatsuba_add2_io_s[193:0]                         ), //o
    .clk    (clk                                                ), //i
    .resetn (resetn                                             )  //i
  );
  BADD_1672 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[287:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[287:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[288:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[192:0];
  assign karatsuba_noExtend_add3_io_a = {95'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[95 : 0] = _zz_io_b;
    karatsuba_noExtend_add3_io_b[287 : 96] = karatsuba_msbMul_karatsuba_msbMul_io_p_delay_5;
  end

  always @(*) begin
    io_p[95 : 0] = _zz_io_p_1;
    io_p[383 : 96] = karatsuba_noExtend_add3_io_s[287:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_a_1 <= karatsuba_midAdd_0_1_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b_1 <= karatsuba_midAdd_1_1_io_S;
    karatsuba_msbMul_karatsuba_add1_io_s_delay_1 <= karatsuba_add1_io_s;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 96);
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_5 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4;
    _zz_io_p <= karatsuba_lsbMul_io_p[95 : 0];
    _zz_io_p_1 <= _zz_io_p;
  end


endmodule

module KaratsubaCore_142 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_a_1,
  input      [48:0]   io_a_2,
  input      [48:0]   io_a_3,
  input      [48:0]   io_b_0,
  input      [48:0]   io_b_1,
  input      [48:0]   io_b_2,
  input      [48:0]   io_b_3,
  output reg [385:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [194:0]  karatsuba_add2_io_a;
  wire       [194:0]  karatsuba_hasExtend_add3_io_a;
  wire       [194:0]  karatsuba_hasExtend_add3_io_b;
  wire       [193:0]  karatsuba_hasExtend_add4_io_a;
  wire       [193:0]  karatsuba_lsbMul_io_p;
  wire       [195:0]  karatsuba_midMul_io_p;
  wire       [193:0]  karatsuba_msbMul_io_p;
  wire       [49:0]   karatsuba_midAdd_0_0_io_S;
  wire       [49:0]   karatsuba_midAdd_0_1_io_S;
  wire       [49:0]   karatsuba_midAdd_1_0_io_S;
  wire       [49:0]   karatsuba_midAdd_1_1_io_S;
  wire       [194:0]  karatsuba_add1_io_s;
  wire       [195:0]  karatsuba_add2_io_s;
  wire       [195:0]  karatsuba_hasExtend_add3_io_s;
  wire       [194:0]  karatsuba_hasExtend_add4_io_s;
  wire       [97:0]   _zz_io_b;
  wire       [99:0]   _zz_io_a;
  reg        [49:0]   _zz_io_a_0;
  reg        [49:0]   _zz_io_a_1;
  reg        [49:0]   _zz_io_b_0;
  reg        [49:0]   _zz_io_b_1;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_4;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_5;
  reg        [95:0]   _zz_io_p;
  reg        [95:0]   _zz_io_p_1;
  reg        [95:0]   _zz_io_p_2;

  assign _zz_io_b = (karatsuba_lsbMul_io_p >>> 96);
  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 96);
  KaratsubaCore_462 karatsuba_lsbMul (
    .io_a_0 (io_a_0[48:0]                ), //i
    .io_a_1 (io_a_1[48:0]                ), //i
    .io_b_0 (io_b_0[48:0]                ), //i
    .io_b_1 (io_b_1[48:0]                ), //i
    .io_p   (karatsuba_lsbMul_io_p[193:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_463 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[49:0]            ), //i
    .io_a_1 (_zz_io_a_1[49:0]            ), //i
    .io_b_0 (_zz_io_b_0[49:0]            ), //i
    .io_b_1 (_zz_io_b_1[49:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[195:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_464 karatsuba_msbMul (
    .io_a_0 (io_a_2[48:0]                ), //i
    .io_a_1 (io_a_3[48:0]                ), //i
    .io_b_0 (io_b_2[48:0]                ), //i
    .io_b_1 (io_b_3[48:0]                ), //i
    .io_p   (karatsuba_msbMul_io_p[193:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  ADD_8288 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[48:0]                   ), //i
    .io_A_1 (io_a_2[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[49:0])  //o
  );
  ADD_8288 karatsuba_midAdd_0_1 (
    .io_A_0 (io_a_1[48:0]                   ), //i
    .io_A_1 (io_a_3[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_1_io_S[49:0])  //o
  );
  ADD_8288 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[48:0]                   ), //i
    .io_A_1 (io_b_2[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[49:0])  //o
  );
  ADD_8288 karatsuba_midAdd_1_1 (
    .io_A_0 (io_b_1[48:0]                   ), //i
    .io_A_1 (io_b_3[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_1_io_S[49:0])  //o
  );
  BADD_1666 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[193:0]), //i
    .io_b   (karatsuba_msbMul_io_p[193:0]), //i
    .io_c   (1'b0                        ), //i
    .io_s   (karatsuba_add1_io_s[194:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_1667 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[194:0]), //i
    .io_b   (karatsuba_add1_io_s[194:0]), //i
    .io_c   (1'b1                      ), //i
    .io_s   (karatsuba_add2_io_s[195:0]), //o
    .clk    (clk                       ), //i
    .resetn (resetn                    )  //i
  );
  BADD_1668 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[194:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[194:0]), //i
    .io_c   (1'b0                                ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[195:0]), //o
    .clk    (clk                                 ), //i
    .resetn (resetn                              )  //i
  );
  BADD_1666 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[193:0]                 ), //i
    .io_b   (karatsuba_midMul_karatsuba_msbMul_io_p_delay_5[193:0]), //i
    .io_c   (1'b0                                                 ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[194:0]                 ), //o
    .clk    (clk                                                  ), //i
    .resetn (resetn                                               )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[194:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[194:0];
  assign karatsuba_hasExtend_add3_io_b = {97'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {94'd0, _zz_io_a};
  always @(*) begin
    io_p[95 : 0] = _zz_io_p_1;
    io_p[191 : 96] = _zz_io_p_2;
    io_p[385 : 192] = karatsuba_hasExtend_add4_io_s[193:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_a_1 <= karatsuba_midAdd_0_1_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b_1 <= karatsuba_midAdd_1_1_io_S;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_5 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_4;
    _zz_io_p <= karatsuba_lsbMul_io_p[95 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= karatsuba_hasExtend_add3_io_s[95:0];
  end


endmodule

module KaratsubaCore_141 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_a_2,
  input      [47:0]   io_a_3,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  input      [47:0]   io_b_2,
  input      [47:0]   io_b_3,
  output reg [383:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [192:0]  karatsuba_add2_io_a;
  wire       [287:0]  karatsuba_noExtend_add3_io_a;
  reg        [287:0]  karatsuba_noExtend_add3_io_b;
  wire       [191:0]  karatsuba_lsbMul_io_p;
  wire       [193:0]  karatsuba_midMul_io_p;
  wire       [191:0]  karatsuba_msbMul_io_p;
  wire       [48:0]   karatsuba_midAdd_0_0_io_S;
  wire       [48:0]   karatsuba_midAdd_0_1_io_S;
  wire       [48:0]   karatsuba_midAdd_1_0_io_S;
  wire       [48:0]   karatsuba_midAdd_1_1_io_S;
  wire       [192:0]  karatsuba_add1_io_s;
  wire       [193:0]  karatsuba_add2_io_s;
  wire       [288:0]  karatsuba_noExtend_add3_io_s;
  wire       [192:0]  _zz_io_a;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_a_1;
  reg        [48:0]   _zz_io_b_0;
  reg        [48:0]   _zz_io_b_1;
  reg        [192:0]  karatsuba_lsbMul_karatsuba_add1_io_s_delay_1;
  reg        [95:0]   _zz_io_b;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_5;
  reg        [95:0]   _zz_io_p;
  reg        [95:0]   _zz_io_p_1;

  assign _zz_io_a = karatsuba_add2_io_s[192:0];
  KaratsubaCore_465 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]                ), //i
    .io_a_1 (io_a_1[47:0]                ), //i
    .io_b_0 (io_b_0[47:0]                ), //i
    .io_b_1 (io_b_1[47:0]                ), //i
    .io_p   (karatsuba_lsbMul_io_p[191:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_466 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]            ), //i
    .io_a_1 (_zz_io_a_1[48:0]            ), //i
    .io_b_0 (_zz_io_b_0[48:0]            ), //i
    .io_b_1 (_zz_io_b_1[48:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[193:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_467 karatsuba_msbMul (
    .io_a_0 (io_a_2[47:0]                ), //i
    .io_a_1 (io_a_3[47:0]                ), //i
    .io_b_0 (io_b_2[47:0]                ), //i
    .io_b_1 (io_b_3[47:0]                ), //i
    .io_p   (karatsuba_msbMul_io_p[191:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  ADD_11602 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[47:0]                   ), //i
    .io_A_1 (io_a_2[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_0_1 (
    .io_A_0 (io_a_1[47:0]                   ), //i
    .io_A_1 (io_a_3[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_1_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[47:0]                   ), //i
    .io_A_1 (io_b_2[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_1 (
    .io_A_0 (io_b_1[47:0]                   ), //i
    .io_A_1 (io_b_3[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_1_io_S[48:0])  //o
  );
  BADD_1670 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[191:0]), //i
    .io_b   (karatsuba_msbMul_io_p[191:0]), //i
    .io_c   (1'b0                        ), //i
    .io_s   (karatsuba_add1_io_s[192:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_1671 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[192:0]                         ), //i
    .io_b   (karatsuba_lsbMul_karatsuba_add1_io_s_delay_1[192:0]), //i
    .io_c   (1'b1                                               ), //i
    .io_s   (karatsuba_add2_io_s[193:0]                         ), //o
    .clk    (clk                                                ), //i
    .resetn (resetn                                             )  //i
  );
  BADD_1672 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[287:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[287:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[288:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[192:0];
  assign karatsuba_noExtend_add3_io_a = {95'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[95 : 0] = _zz_io_b;
    karatsuba_noExtend_add3_io_b[287 : 96] = karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_5;
  end

  always @(*) begin
    io_p[95 : 0] = _zz_io_p_1;
    io_p[383 : 96] = karatsuba_noExtend_add3_io_s[287:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_a_1 <= karatsuba_midAdd_0_1_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b_1 <= karatsuba_midAdd_1_1_io_S;
    karatsuba_lsbMul_karatsuba_add1_io_s_delay_1 <= karatsuba_add1_io_s;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 96);
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_5 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4;
    _zz_io_p <= karatsuba_lsbMul_io_p[95 : 0];
    _zz_io_p_1 <= _zz_io_p;
  end


endmodule

//ADD_4265 replaced by ADD_5761

//ADD_4264 replaced by ADD_5756

//ADD_4263 replaced by ADD_5756

//ADD_4262 replaced by ADD_5756

//ADD_4261 replaced by ADD_5756

//ADD_4260 replaced by ADD_5756

//ADD_4277 replaced by ADD_11602

//ADD_4276 replaced by ADD_11602

//ADD_4275 replaced by ADD_11602

//ADD_4274 replaced by ADD_11602

//ADD_4273 replaced by ADD_11602

//ADD_4272 replaced by ADD_11602

//ADD_4271 replaced by ADD_11602

//ADD_4270 replaced by ADD_11602

//ADD_4269 replaced by ADD_11602

//ADD_4268 replaced by ADD_11602

//ADD_4267 replaced by ADD_11602

//ADD_4266 replaced by ADD_11602

//ADD_4286 replaced by ADD_11601

//ADD_4285 replaced by ADD_11602

//ADD_4284 replaced by ADD_11602

//ADD_4283 replaced by ADD_11602

//ADD_4282 replaced by ADD_11602

//ADD_4281 replaced by ADD_11602

//ADD_4280 replaced by ADD_11602

//ADD_4279 replaced by ADD_11602

//ADD_4278 replaced by ADD_11602

//ADD_4294 replaced by ADD_11602

//ADD_4293 replaced by ADD_11602

//ADD_4292 replaced by ADD_11602

//ADD_4291 replaced by ADD_11602

//ADD_4290 replaced by ADD_11602

//ADD_4289 replaced by ADD_11602

//ADD_4288 replaced by ADD_11602

//ADD_4287 replaced by ADD_11602

//BADD_1315 replaced by BADD_1672

//BADD_1314 replaced by BADD_1671

//BADD_1313 replaced by BADD_1670

//ADD_4298 replaced by ADD_11602

//ADD_4297 replaced by ADD_11602

//ADD_4296 replaced by ADD_11602

//ADD_4295 replaced by ADD_11602

//KaratsubaCore_146 replaced by KaratsubaCore_467

//KaratsubaCore_145 replaced by KaratsubaCore_466

//KaratsubaCore_144 replaced by KaratsubaCore_465

//BADD_1319 replaced by BADD_1666

//BADD_1318 replaced by BADD_1668

//BADD_1317 replaced by BADD_1667

//BADD_1316 replaced by BADD_1666

//ADD_4302 replaced by ADD_8288

//ADD_4301 replaced by ADD_8288

//ADD_4300 replaced by ADD_8288

//ADD_4299 replaced by ADD_8288

//KaratsubaCore_149 replaced by KaratsubaCore_464

//KaratsubaCore_148 replaced by KaratsubaCore_463

//KaratsubaCore_147 replaced by KaratsubaCore_462

//BADD_1322 replaced by BADD_1672

//BADD_1321 replaced by BADD_1671

//BADD_1320 replaced by BADD_1670

//ADD_4306 replaced by ADD_11602

//ADD_4305 replaced by ADD_11602

//ADD_4304 replaced by ADD_11602

//ADD_4303 replaced by ADD_11602

//KaratsubaCore_152 replaced by KaratsubaCore_467

//KaratsubaCore_151 replaced by KaratsubaCore_466

//KaratsubaCore_150 replaced by KaratsubaCore_465

//ADD_4318 replaced by ADD_11602

//ADD_4317 replaced by ADD_11602

//ADD_4316 replaced by ADD_11602

//ADD_4315 replaced by ADD_11602

//ADD_4314 replaced by ADD_11602

//ADD_4313 replaced by ADD_11602

//ADD_4312 replaced by ADD_11602

//ADD_4311 replaced by ADD_11602

//ADD_4310 replaced by ADD_11602

//ADD_4309 replaced by ADD_11602

//ADD_4308 replaced by ADD_11602

//ADD_4307 replaced by ADD_11602

//ADD_4327 replaced by ADD_11601

//ADD_4326 replaced by ADD_11602

//ADD_4325 replaced by ADD_11602

//ADD_4324 replaced by ADD_11602

//ADD_4323 replaced by ADD_11602

//ADD_4322 replaced by ADD_11602

//ADD_4321 replaced by ADD_11602

//ADD_4320 replaced by ADD_11602

//ADD_4319 replaced by ADD_11602

//ADD_4335 replaced by ADD_11602

//ADD_4334 replaced by ADD_11602

//ADD_4333 replaced by ADD_11602

//ADD_4332 replaced by ADD_11602

//ADD_4331 replaced by ADD_11602

//ADD_4330 replaced by ADD_11602

//ADD_4329 replaced by ADD_11602

//ADD_4328 replaced by ADD_11602

//BADD_1325 replaced by BADD_1672

//BADD_1324 replaced by BADD_1671

//BADD_1323 replaced by BADD_1670

//ADD_4339 replaced by ADD_11602

//ADD_4338 replaced by ADD_11602

//ADD_4337 replaced by ADD_11602

//ADD_4336 replaced by ADD_11602

//KaratsubaCore_155 replaced by KaratsubaCore_467

//KaratsubaCore_154 replaced by KaratsubaCore_466

//KaratsubaCore_153 replaced by KaratsubaCore_465

//BADD_1329 replaced by BADD_1666

//BADD_1328 replaced by BADD_1668

//BADD_1327 replaced by BADD_1667

//BADD_1326 replaced by BADD_1666

//ADD_4343 replaced by ADD_8288

//ADD_4342 replaced by ADD_8288

//ADD_4341 replaced by ADD_8288

//ADD_4340 replaced by ADD_8288

//KaratsubaCore_158 replaced by KaratsubaCore_464

//KaratsubaCore_157 replaced by KaratsubaCore_463

//KaratsubaCore_156 replaced by KaratsubaCore_462

//BADD_1332 replaced by BADD_1672

//BADD_1331 replaced by BADD_1671

//BADD_1330 replaced by BADD_1670

//ADD_4347 replaced by ADD_11602

//ADD_4346 replaced by ADD_11602

//ADD_4345 replaced by ADD_11602

//ADD_4344 replaced by ADD_11602

//KaratsubaCore_161 replaced by KaratsubaCore_467

//KaratsubaCore_160 replaced by KaratsubaCore_466

//KaratsubaCore_159 replaced by KaratsubaCore_465

//ADD_4353 replaced by ADD_5761

//ADD_4352 replaced by ADD_5756

//ADD_4351 replaced by ADD_5756

//ADD_4350 replaced by ADD_5756

//ADD_4349 replaced by ADD_5756

//ADD_4348 replaced by ADD_5756

//ADD_4365 replaced by ADD_11602

//ADD_4364 replaced by ADD_11602

//ADD_4363 replaced by ADD_11602

//ADD_4362 replaced by ADD_11602

//ADD_4361 replaced by ADD_11602

//ADD_4360 replaced by ADD_11602

//ADD_4359 replaced by ADD_11602

//ADD_4358 replaced by ADD_11602

//ADD_4357 replaced by ADD_11602

//ADD_4356 replaced by ADD_11602

//ADD_4355 replaced by ADD_11602

//ADD_4354 replaced by ADD_11602

//ADD_4374 replaced by ADD_11601

//ADD_4373 replaced by ADD_11602

//ADD_4372 replaced by ADD_11602

//ADD_4371 replaced by ADD_11602

//ADD_4370 replaced by ADD_11602

//ADD_4369 replaced by ADD_11602

//ADD_4368 replaced by ADD_11602

//ADD_4367 replaced by ADD_11602

//ADD_4366 replaced by ADD_11602

//ADD_4382 replaced by ADD_11602

//ADD_4381 replaced by ADD_11602

//ADD_4380 replaced by ADD_11602

//ADD_4379 replaced by ADD_11602

//ADD_4378 replaced by ADD_11602

//ADD_4377 replaced by ADD_11602

//ADD_4376 replaced by ADD_11602

//ADD_4375 replaced by ADD_11602

//BADD_1335 replaced by BADD_1672

//BADD_1334 replaced by BADD_1671

//BADD_1333 replaced by BADD_1670

//ADD_4386 replaced by ADD_11602

//ADD_4385 replaced by ADD_11602

//ADD_4384 replaced by ADD_11602

//ADD_4383 replaced by ADD_11602

//KaratsubaCore_164 replaced by KaratsubaCore_467

//KaratsubaCore_163 replaced by KaratsubaCore_466

//KaratsubaCore_162 replaced by KaratsubaCore_465

//BADD_1339 replaced by BADD_1666

//BADD_1338 replaced by BADD_1668

//BADD_1337 replaced by BADD_1667

//BADD_1336 replaced by BADD_1666

//ADD_4390 replaced by ADD_8288

//ADD_4389 replaced by ADD_8288

//ADD_4388 replaced by ADD_8288

//ADD_4387 replaced by ADD_8288

//KaratsubaCore_167 replaced by KaratsubaCore_464

//KaratsubaCore_166 replaced by KaratsubaCore_463

//KaratsubaCore_165 replaced by KaratsubaCore_462

//BADD_1342 replaced by BADD_1672

//BADD_1341 replaced by BADD_1671

//BADD_1340 replaced by BADD_1670

//ADD_4394 replaced by ADD_11602

//ADD_4393 replaced by ADD_11602

//ADD_4392 replaced by ADD_11602

//ADD_4391 replaced by ADD_11602

//KaratsubaCore_170 replaced by KaratsubaCore_467

//KaratsubaCore_169 replaced by KaratsubaCore_466

//KaratsubaCore_168 replaced by KaratsubaCore_465

//ADD_4406 replaced by ADD_11602

//ADD_4405 replaced by ADD_11602

//ADD_4404 replaced by ADD_11602

//ADD_4403 replaced by ADD_11602

//ADD_4402 replaced by ADD_11602

//ADD_4401 replaced by ADD_11602

//ADD_4400 replaced by ADD_11602

//ADD_4399 replaced by ADD_11602

//ADD_4398 replaced by ADD_11602

//ADD_4397 replaced by ADD_11602

//ADD_4396 replaced by ADD_11602

//ADD_4395 replaced by ADD_11602

//ADD_4415 replaced by ADD_11601

//ADD_4414 replaced by ADD_11602

//ADD_4413 replaced by ADD_11602

//ADD_4412 replaced by ADD_11602

//ADD_4411 replaced by ADD_11602

//ADD_4410 replaced by ADD_11602

//ADD_4409 replaced by ADD_11602

//ADD_4408 replaced by ADD_11602

//ADD_4407 replaced by ADD_11602

//ADD_4423 replaced by ADD_11602

//ADD_4422 replaced by ADD_11602

//ADD_4421 replaced by ADD_11602

//ADD_4420 replaced by ADD_11602

//ADD_4419 replaced by ADD_11602

//ADD_4418 replaced by ADD_11602

//ADD_4417 replaced by ADD_11602

//ADD_4416 replaced by ADD_11602

//BADD_1345 replaced by BADD_1672

//BADD_1344 replaced by BADD_1671

//BADD_1343 replaced by BADD_1670

//ADD_4427 replaced by ADD_11602

//ADD_4426 replaced by ADD_11602

//ADD_4425 replaced by ADD_11602

//ADD_4424 replaced by ADD_11602

//KaratsubaCore_173 replaced by KaratsubaCore_467

//KaratsubaCore_172 replaced by KaratsubaCore_466

//KaratsubaCore_171 replaced by KaratsubaCore_465

//BADD_1349 replaced by BADD_1666

//BADD_1348 replaced by BADD_1668

//BADD_1347 replaced by BADD_1667

//BADD_1346 replaced by BADD_1666

//ADD_4431 replaced by ADD_8288

//ADD_4430 replaced by ADD_8288

//ADD_4429 replaced by ADD_8288

//ADD_4428 replaced by ADD_8288

//KaratsubaCore_176 replaced by KaratsubaCore_464

//KaratsubaCore_175 replaced by KaratsubaCore_463

//KaratsubaCore_174 replaced by KaratsubaCore_462

//BADD_1352 replaced by BADD_1672

//BADD_1351 replaced by BADD_1671

//BADD_1350 replaced by BADD_1670

//ADD_4435 replaced by ADD_11602

//ADD_4434 replaced by ADD_11602

//ADD_4433 replaced by ADD_11602

//ADD_4432 replaced by ADD_11602

//KaratsubaCore_179 replaced by KaratsubaCore_467

//KaratsubaCore_178 replaced by KaratsubaCore_466

//KaratsubaCore_177 replaced by KaratsubaCore_465

//ADD_4441 replaced by ADD_5761

//ADD_4440 replaced by ADD_5756

//ADD_4439 replaced by ADD_5756

//ADD_4438 replaced by ADD_5756

//ADD_4437 replaced by ADD_5756

//ADD_4436 replaced by ADD_5756

//ADD_4453 replaced by ADD_11602

//ADD_4452 replaced by ADD_11602

//ADD_4451 replaced by ADD_11602

//ADD_4450 replaced by ADD_11602

//ADD_4449 replaced by ADD_11602

//ADD_4448 replaced by ADD_11602

//ADD_4447 replaced by ADD_11602

//ADD_4446 replaced by ADD_11602

//ADD_4445 replaced by ADD_11602

//ADD_4444 replaced by ADD_11602

//ADD_4443 replaced by ADD_11602

//ADD_4442 replaced by ADD_11602

//ADD_4462 replaced by ADD_11601

//ADD_4461 replaced by ADD_11602

//ADD_4460 replaced by ADD_11602

//ADD_4459 replaced by ADD_11602

//ADD_4458 replaced by ADD_11602

//ADD_4457 replaced by ADD_11602

//ADD_4456 replaced by ADD_11602

//ADD_4455 replaced by ADD_11602

//ADD_4454 replaced by ADD_11602

//ADD_4470 replaced by ADD_11602

//ADD_4469 replaced by ADD_11602

//ADD_4468 replaced by ADD_11602

//ADD_4467 replaced by ADD_11602

//ADD_4466 replaced by ADD_11602

//ADD_4465 replaced by ADD_11602

//ADD_4464 replaced by ADD_11602

//ADD_4463 replaced by ADD_11602

//BADD_1355 replaced by BADD_1672

//BADD_1354 replaced by BADD_1671

//BADD_1353 replaced by BADD_1670

//ADD_4474 replaced by ADD_11602

//ADD_4473 replaced by ADD_11602

//ADD_4472 replaced by ADD_11602

//ADD_4471 replaced by ADD_11602

//KaratsubaCore_182 replaced by KaratsubaCore_467

//KaratsubaCore_181 replaced by KaratsubaCore_466

//KaratsubaCore_180 replaced by KaratsubaCore_465

//BADD_1359 replaced by BADD_1666

//BADD_1358 replaced by BADD_1668

//BADD_1357 replaced by BADD_1667

//BADD_1356 replaced by BADD_1666

//ADD_4478 replaced by ADD_8288

//ADD_4477 replaced by ADD_8288

//ADD_4476 replaced by ADD_8288

//ADD_4475 replaced by ADD_8288

//KaratsubaCore_185 replaced by KaratsubaCore_464

//KaratsubaCore_184 replaced by KaratsubaCore_463

//KaratsubaCore_183 replaced by KaratsubaCore_462

//BADD_1362 replaced by BADD_1672

//BADD_1361 replaced by BADD_1671

//BADD_1360 replaced by BADD_1670

//ADD_4482 replaced by ADD_11602

//ADD_4481 replaced by ADD_11602

//ADD_4480 replaced by ADD_11602

//ADD_4479 replaced by ADD_11602

//KaratsubaCore_188 replaced by KaratsubaCore_467

//KaratsubaCore_187 replaced by KaratsubaCore_466

//KaratsubaCore_186 replaced by KaratsubaCore_465

//ADD_4494 replaced by ADD_11602

//ADD_4493 replaced by ADD_11602

//ADD_4492 replaced by ADD_11602

//ADD_4491 replaced by ADD_11602

//ADD_4490 replaced by ADD_11602

//ADD_4489 replaced by ADD_11602

//ADD_4488 replaced by ADD_11602

//ADD_4487 replaced by ADD_11602

//ADD_4486 replaced by ADD_11602

//ADD_4485 replaced by ADD_11602

//ADD_4484 replaced by ADD_11602

//ADD_4483 replaced by ADD_11602

//ADD_4503 replaced by ADD_11601

//ADD_4502 replaced by ADD_11602

//ADD_4501 replaced by ADD_11602

//ADD_4500 replaced by ADD_11602

//ADD_4499 replaced by ADD_11602

//ADD_4498 replaced by ADD_11602

//ADD_4497 replaced by ADD_11602

//ADD_4496 replaced by ADD_11602

//ADD_4495 replaced by ADD_11602

//ADD_4511 replaced by ADD_11602

//ADD_4510 replaced by ADD_11602

//ADD_4509 replaced by ADD_11602

//ADD_4508 replaced by ADD_11602

//ADD_4507 replaced by ADD_11602

//ADD_4506 replaced by ADD_11602

//ADD_4505 replaced by ADD_11602

//ADD_4504 replaced by ADD_11602

//BADD_1365 replaced by BADD_1672

//BADD_1364 replaced by BADD_1671

//BADD_1363 replaced by BADD_1670

//ADD_4515 replaced by ADD_11602

//ADD_4514 replaced by ADD_11602

//ADD_4513 replaced by ADD_11602

//ADD_4512 replaced by ADD_11602

//KaratsubaCore_191 replaced by KaratsubaCore_467

//KaratsubaCore_190 replaced by KaratsubaCore_466

//KaratsubaCore_189 replaced by KaratsubaCore_465

//BADD_1369 replaced by BADD_1666

//BADD_1368 replaced by BADD_1668

//BADD_1367 replaced by BADD_1667

//BADD_1366 replaced by BADD_1666

//ADD_4519 replaced by ADD_8288

//ADD_4518 replaced by ADD_8288

//ADD_4517 replaced by ADD_8288

//ADD_4516 replaced by ADD_8288

//KaratsubaCore_194 replaced by KaratsubaCore_464

//KaratsubaCore_193 replaced by KaratsubaCore_463

//KaratsubaCore_192 replaced by KaratsubaCore_462

//BADD_1372 replaced by BADD_1672

//BADD_1371 replaced by BADD_1671

//BADD_1370 replaced by BADD_1670

//ADD_4523 replaced by ADD_11602

//ADD_4522 replaced by ADD_11602

//ADD_4521 replaced by ADD_11602

//ADD_4520 replaced by ADD_11602

//KaratsubaCore_197 replaced by KaratsubaCore_467

//KaratsubaCore_196 replaced by KaratsubaCore_466

//KaratsubaCore_195 replaced by KaratsubaCore_465

//ADD_4529 replaced by ADD_5761

//ADD_4528 replaced by ADD_5756

//ADD_4527 replaced by ADD_5756

//ADD_4526 replaced by ADD_5756

//ADD_4525 replaced by ADD_5756

//ADD_4524 replaced by ADD_5756

//ADD_4541 replaced by ADD_11602

//ADD_4540 replaced by ADD_11602

//ADD_4539 replaced by ADD_11602

//ADD_4538 replaced by ADD_11602

//ADD_4537 replaced by ADD_11602

//ADD_4536 replaced by ADD_11602

//ADD_4535 replaced by ADD_11602

//ADD_4534 replaced by ADD_11602

//ADD_4533 replaced by ADD_11602

//ADD_4532 replaced by ADD_11602

//ADD_4531 replaced by ADD_11602

//ADD_4530 replaced by ADD_11602

//ADD_4550 replaced by ADD_11601

//ADD_4549 replaced by ADD_11602

//ADD_4548 replaced by ADD_11602

//ADD_4547 replaced by ADD_11602

//ADD_4546 replaced by ADD_11602

//ADD_4545 replaced by ADD_11602

//ADD_4544 replaced by ADD_11602

//ADD_4543 replaced by ADD_11602

//ADD_4542 replaced by ADD_11602

//ADD_4558 replaced by ADD_11602

//ADD_4557 replaced by ADD_11602

//ADD_4556 replaced by ADD_11602

//ADD_4555 replaced by ADD_11602

//ADD_4554 replaced by ADD_11602

//ADD_4553 replaced by ADD_11602

//ADD_4552 replaced by ADD_11602

//ADD_4551 replaced by ADD_11602

//BADD_1375 replaced by BADD_1672

//BADD_1374 replaced by BADD_1671

//BADD_1373 replaced by BADD_1670

//ADD_4562 replaced by ADD_11602

//ADD_4561 replaced by ADD_11602

//ADD_4560 replaced by ADD_11602

//ADD_4559 replaced by ADD_11602

//KaratsubaCore_200 replaced by KaratsubaCore_467

//KaratsubaCore_199 replaced by KaratsubaCore_466

//KaratsubaCore_198 replaced by KaratsubaCore_465

//BADD_1379 replaced by BADD_1666

//BADD_1378 replaced by BADD_1668

//BADD_1377 replaced by BADD_1667

//BADD_1376 replaced by BADD_1666

//ADD_4566 replaced by ADD_8288

//ADD_4565 replaced by ADD_8288

//ADD_4564 replaced by ADD_8288

//ADD_4563 replaced by ADD_8288

//KaratsubaCore_203 replaced by KaratsubaCore_464

//KaratsubaCore_202 replaced by KaratsubaCore_463

//KaratsubaCore_201 replaced by KaratsubaCore_462

//BADD_1382 replaced by BADD_1672

//BADD_1381 replaced by BADD_1671

//BADD_1380 replaced by BADD_1670

//ADD_4570 replaced by ADD_11602

//ADD_4569 replaced by ADD_11602

//ADD_4568 replaced by ADD_11602

//ADD_4567 replaced by ADD_11602

//KaratsubaCore_206 replaced by KaratsubaCore_467

//KaratsubaCore_205 replaced by KaratsubaCore_466

//KaratsubaCore_204 replaced by KaratsubaCore_465

//ADD_4582 replaced by ADD_11602

//ADD_4581 replaced by ADD_11602

//ADD_4580 replaced by ADD_11602

//ADD_4579 replaced by ADD_11602

//ADD_4578 replaced by ADD_11602

//ADD_4577 replaced by ADD_11602

//ADD_4576 replaced by ADD_11602

//ADD_4575 replaced by ADD_11602

//ADD_4574 replaced by ADD_11602

//ADD_4573 replaced by ADD_11602

//ADD_4572 replaced by ADD_11602

//ADD_4571 replaced by ADD_11602

//ADD_4591 replaced by ADD_11601

//ADD_4590 replaced by ADD_11602

//ADD_4589 replaced by ADD_11602

//ADD_4588 replaced by ADD_11602

//ADD_4587 replaced by ADD_11602

//ADD_4586 replaced by ADD_11602

//ADD_4585 replaced by ADD_11602

//ADD_4584 replaced by ADD_11602

//ADD_4583 replaced by ADD_11602

//ADD_4599 replaced by ADD_11602

//ADD_4598 replaced by ADD_11602

//ADD_4597 replaced by ADD_11602

//ADD_4596 replaced by ADD_11602

//ADD_4595 replaced by ADD_11602

//ADD_4594 replaced by ADD_11602

//ADD_4593 replaced by ADD_11602

//ADD_4592 replaced by ADD_11602

//BADD_1385 replaced by BADD_1672

//BADD_1384 replaced by BADD_1671

//BADD_1383 replaced by BADD_1670

//ADD_4603 replaced by ADD_11602

//ADD_4602 replaced by ADD_11602

//ADD_4601 replaced by ADD_11602

//ADD_4600 replaced by ADD_11602

//KaratsubaCore_209 replaced by KaratsubaCore_467

//KaratsubaCore_208 replaced by KaratsubaCore_466

//KaratsubaCore_207 replaced by KaratsubaCore_465

//BADD_1389 replaced by BADD_1666

//BADD_1388 replaced by BADD_1668

//BADD_1387 replaced by BADD_1667

//BADD_1386 replaced by BADD_1666

//ADD_4607 replaced by ADD_8288

//ADD_4606 replaced by ADD_8288

//ADD_4605 replaced by ADD_8288

//ADD_4604 replaced by ADD_8288

//KaratsubaCore_212 replaced by KaratsubaCore_464

//KaratsubaCore_211 replaced by KaratsubaCore_463

//KaratsubaCore_210 replaced by KaratsubaCore_462

//BADD_1392 replaced by BADD_1672

//BADD_1391 replaced by BADD_1671

//BADD_1390 replaced by BADD_1670

//ADD_4611 replaced by ADD_11602

//ADD_4610 replaced by ADD_11602

//ADD_4609 replaced by ADD_11602

//ADD_4608 replaced by ADD_11602

//KaratsubaCore_215 replaced by KaratsubaCore_467

//KaratsubaCore_214 replaced by KaratsubaCore_466

//KaratsubaCore_213 replaced by KaratsubaCore_465

//ADD_4617 replaced by ADD_5761

//ADD_4616 replaced by ADD_5756

//ADD_4615 replaced by ADD_5756

//ADD_4614 replaced by ADD_5756

//ADD_4613 replaced by ADD_5756

//ADD_4612 replaced by ADD_5756

//ADD_4629 replaced by ADD_11602

//ADD_4628 replaced by ADD_11602

//ADD_4627 replaced by ADD_11602

//ADD_4626 replaced by ADD_11602

//ADD_4625 replaced by ADD_11602

//ADD_4624 replaced by ADD_11602

//ADD_4623 replaced by ADD_11602

//ADD_4622 replaced by ADD_11602

//ADD_4621 replaced by ADD_11602

//ADD_4620 replaced by ADD_11602

//ADD_4619 replaced by ADD_11602

//ADD_4618 replaced by ADD_11602

//ADD_4638 replaced by ADD_11601

//ADD_4637 replaced by ADD_11602

//ADD_4636 replaced by ADD_11602

//ADD_4635 replaced by ADD_11602

//ADD_4634 replaced by ADD_11602

//ADD_4633 replaced by ADD_11602

//ADD_4632 replaced by ADD_11602

//ADD_4631 replaced by ADD_11602

//ADD_4630 replaced by ADD_11602

//ADD_4646 replaced by ADD_11602

//ADD_4645 replaced by ADD_11602

//ADD_4644 replaced by ADD_11602

//ADD_4643 replaced by ADD_11602

//ADD_4642 replaced by ADD_11602

//ADD_4641 replaced by ADD_11602

//ADD_4640 replaced by ADD_11602

//ADD_4639 replaced by ADD_11602

//BADD_1395 replaced by BADD_1672

//BADD_1394 replaced by BADD_1671

//BADD_1393 replaced by BADD_1670

//ADD_4650 replaced by ADD_11602

//ADD_4649 replaced by ADD_11602

//ADD_4648 replaced by ADD_11602

//ADD_4647 replaced by ADD_11602

//KaratsubaCore_218 replaced by KaratsubaCore_467

//KaratsubaCore_217 replaced by KaratsubaCore_466

//KaratsubaCore_216 replaced by KaratsubaCore_465

//BADD_1399 replaced by BADD_1666

//BADD_1398 replaced by BADD_1668

//BADD_1397 replaced by BADD_1667

//BADD_1396 replaced by BADD_1666

//ADD_4654 replaced by ADD_8288

//ADD_4653 replaced by ADD_8288

//ADD_4652 replaced by ADD_8288

//ADD_4651 replaced by ADD_8288

//KaratsubaCore_221 replaced by KaratsubaCore_464

//KaratsubaCore_220 replaced by KaratsubaCore_463

//KaratsubaCore_219 replaced by KaratsubaCore_462

//BADD_1402 replaced by BADD_1672

//BADD_1401 replaced by BADD_1671

//BADD_1400 replaced by BADD_1670

//ADD_4658 replaced by ADD_11602

//ADD_4657 replaced by ADD_11602

//ADD_4656 replaced by ADD_11602

//ADD_4655 replaced by ADD_11602

//KaratsubaCore_224 replaced by KaratsubaCore_467

//KaratsubaCore_223 replaced by KaratsubaCore_466

//KaratsubaCore_222 replaced by KaratsubaCore_465

//ADD_4670 replaced by ADD_11602

//ADD_4669 replaced by ADD_11602

//ADD_4668 replaced by ADD_11602

//ADD_4667 replaced by ADD_11602

//ADD_4666 replaced by ADD_11602

//ADD_4665 replaced by ADD_11602

//ADD_4664 replaced by ADD_11602

//ADD_4663 replaced by ADD_11602

//ADD_4662 replaced by ADD_11602

//ADD_4661 replaced by ADD_11602

//ADD_4660 replaced by ADD_11602

//ADD_4659 replaced by ADD_11602

//ADD_4679 replaced by ADD_11601

//ADD_4678 replaced by ADD_11602

//ADD_4677 replaced by ADD_11602

//ADD_4676 replaced by ADD_11602

//ADD_4675 replaced by ADD_11602

//ADD_4674 replaced by ADD_11602

//ADD_4673 replaced by ADD_11602

//ADD_4672 replaced by ADD_11602

//ADD_4671 replaced by ADD_11602

//ADD_4687 replaced by ADD_11602

//ADD_4686 replaced by ADD_11602

//ADD_4685 replaced by ADD_11602

//ADD_4684 replaced by ADD_11602

//ADD_4683 replaced by ADD_11602

//ADD_4682 replaced by ADD_11602

//ADD_4681 replaced by ADD_11602

//ADD_4680 replaced by ADD_11602

//BADD_1405 replaced by BADD_1672

//BADD_1404 replaced by BADD_1671

//BADD_1403 replaced by BADD_1670

//ADD_4691 replaced by ADD_11602

//ADD_4690 replaced by ADD_11602

//ADD_4689 replaced by ADD_11602

//ADD_4688 replaced by ADD_11602

//KaratsubaCore_227 replaced by KaratsubaCore_467

//KaratsubaCore_226 replaced by KaratsubaCore_466

//KaratsubaCore_225 replaced by KaratsubaCore_465

//BADD_1409 replaced by BADD_1666

//BADD_1408 replaced by BADD_1668

//BADD_1407 replaced by BADD_1667

//BADD_1406 replaced by BADD_1666

//ADD_4695 replaced by ADD_8288

//ADD_4694 replaced by ADD_8288

//ADD_4693 replaced by ADD_8288

//ADD_4692 replaced by ADD_8288

//KaratsubaCore_230 replaced by KaratsubaCore_464

//KaratsubaCore_229 replaced by KaratsubaCore_463

//KaratsubaCore_228 replaced by KaratsubaCore_462

//BADD_1412 replaced by BADD_1672

//BADD_1411 replaced by BADD_1671

//BADD_1410 replaced by BADD_1670

//ADD_4699 replaced by ADD_11602

//ADD_4698 replaced by ADD_11602

//ADD_4697 replaced by ADD_11602

//ADD_4696 replaced by ADD_11602

//KaratsubaCore_233 replaced by KaratsubaCore_467

//KaratsubaCore_232 replaced by KaratsubaCore_466

//KaratsubaCore_231 replaced by KaratsubaCore_465

//ADD_4705 replaced by ADD_5761

//ADD_4704 replaced by ADD_5756

//ADD_4703 replaced by ADD_5756

//ADD_4702 replaced by ADD_5756

//ADD_4701 replaced by ADD_5756

//ADD_4700 replaced by ADD_5756

//ADD_4717 replaced by ADD_11602

//ADD_4716 replaced by ADD_11602

//ADD_4715 replaced by ADD_11602

//ADD_4714 replaced by ADD_11602

//ADD_4713 replaced by ADD_11602

//ADD_4712 replaced by ADD_11602

//ADD_4711 replaced by ADD_11602

//ADD_4710 replaced by ADD_11602

//ADD_4709 replaced by ADD_11602

//ADD_4708 replaced by ADD_11602

//ADD_4707 replaced by ADD_11602

//ADD_4706 replaced by ADD_11602

//ADD_4726 replaced by ADD_11601

//ADD_4725 replaced by ADD_11602

//ADD_4724 replaced by ADD_11602

//ADD_4723 replaced by ADD_11602

//ADD_4722 replaced by ADD_11602

//ADD_4721 replaced by ADD_11602

//ADD_4720 replaced by ADD_11602

//ADD_4719 replaced by ADD_11602

//ADD_4718 replaced by ADD_11602

//ADD_4734 replaced by ADD_11602

//ADD_4733 replaced by ADD_11602

//ADD_4732 replaced by ADD_11602

//ADD_4731 replaced by ADD_11602

//ADD_4730 replaced by ADD_11602

//ADD_4729 replaced by ADD_11602

//ADD_4728 replaced by ADD_11602

//ADD_4727 replaced by ADD_11602

//BADD_1415 replaced by BADD_1672

//BADD_1414 replaced by BADD_1671

//BADD_1413 replaced by BADD_1670

//ADD_4738 replaced by ADD_11602

//ADD_4737 replaced by ADD_11602

//ADD_4736 replaced by ADD_11602

//ADD_4735 replaced by ADD_11602

//KaratsubaCore_236 replaced by KaratsubaCore_467

//KaratsubaCore_235 replaced by KaratsubaCore_466

//KaratsubaCore_234 replaced by KaratsubaCore_465

//BADD_1419 replaced by BADD_1666

//BADD_1418 replaced by BADD_1668

//BADD_1417 replaced by BADD_1667

//BADD_1416 replaced by BADD_1666

//ADD_4742 replaced by ADD_8288

//ADD_4741 replaced by ADD_8288

//ADD_4740 replaced by ADD_8288

//ADD_4739 replaced by ADD_8288

//KaratsubaCore_239 replaced by KaratsubaCore_464

//KaratsubaCore_238 replaced by KaratsubaCore_463

//KaratsubaCore_237 replaced by KaratsubaCore_462

//BADD_1422 replaced by BADD_1672

//BADD_1421 replaced by BADD_1671

//BADD_1420 replaced by BADD_1670

//ADD_4746 replaced by ADD_11602

//ADD_4745 replaced by ADD_11602

//ADD_4744 replaced by ADD_11602

//ADD_4743 replaced by ADD_11602

//KaratsubaCore_242 replaced by KaratsubaCore_467

//KaratsubaCore_241 replaced by KaratsubaCore_466

//KaratsubaCore_240 replaced by KaratsubaCore_465

//ADD_4758 replaced by ADD_11602

//ADD_4757 replaced by ADD_11602

//ADD_4756 replaced by ADD_11602

//ADD_4755 replaced by ADD_11602

//ADD_4754 replaced by ADD_11602

//ADD_4753 replaced by ADD_11602

//ADD_4752 replaced by ADD_11602

//ADD_4751 replaced by ADD_11602

//ADD_4750 replaced by ADD_11602

//ADD_4749 replaced by ADD_11602

//ADD_4748 replaced by ADD_11602

//ADD_4747 replaced by ADD_11602

//ADD_4767 replaced by ADD_11601

//ADD_4766 replaced by ADD_11602

//ADD_4765 replaced by ADD_11602

//ADD_4764 replaced by ADD_11602

//ADD_4763 replaced by ADD_11602

//ADD_4762 replaced by ADD_11602

//ADD_4761 replaced by ADD_11602

//ADD_4760 replaced by ADD_11602

//ADD_4759 replaced by ADD_11602

//ADD_4775 replaced by ADD_11602

//ADD_4774 replaced by ADD_11602

//ADD_4773 replaced by ADD_11602

//ADD_4772 replaced by ADD_11602

//ADD_4771 replaced by ADD_11602

//ADD_4770 replaced by ADD_11602

//ADD_4769 replaced by ADD_11602

//ADD_4768 replaced by ADD_11602

//BADD_1425 replaced by BADD_1672

//BADD_1424 replaced by BADD_1671

//BADD_1423 replaced by BADD_1670

//ADD_4779 replaced by ADD_11602

//ADD_4778 replaced by ADD_11602

//ADD_4777 replaced by ADD_11602

//ADD_4776 replaced by ADD_11602

//KaratsubaCore_245 replaced by KaratsubaCore_467

//KaratsubaCore_244 replaced by KaratsubaCore_466

//KaratsubaCore_243 replaced by KaratsubaCore_465

//BADD_1429 replaced by BADD_1666

//BADD_1428 replaced by BADD_1668

//BADD_1427 replaced by BADD_1667

//BADD_1426 replaced by BADD_1666

//ADD_4783 replaced by ADD_8288

//ADD_4782 replaced by ADD_8288

//ADD_4781 replaced by ADD_8288

//ADD_4780 replaced by ADD_8288

//KaratsubaCore_248 replaced by KaratsubaCore_464

//KaratsubaCore_247 replaced by KaratsubaCore_463

//KaratsubaCore_246 replaced by KaratsubaCore_462

//BADD_1432 replaced by BADD_1672

//BADD_1431 replaced by BADD_1671

//BADD_1430 replaced by BADD_1670

//ADD_4787 replaced by ADD_11602

//ADD_4786 replaced by ADD_11602

//ADD_4785 replaced by ADD_11602

//ADD_4784 replaced by ADD_11602

//KaratsubaCore_251 replaced by KaratsubaCore_467

//KaratsubaCore_250 replaced by KaratsubaCore_466

//KaratsubaCore_249 replaced by KaratsubaCore_465

//ADD_4793 replaced by ADD_5761

//ADD_4792 replaced by ADD_5756

//ADD_4791 replaced by ADD_5756

//ADD_4790 replaced by ADD_5756

//ADD_4789 replaced by ADD_5756

//ADD_4788 replaced by ADD_5756

//ADD_4805 replaced by ADD_11602

//ADD_4804 replaced by ADD_11602

//ADD_4803 replaced by ADD_11602

//ADD_4802 replaced by ADD_11602

//ADD_4801 replaced by ADD_11602

//ADD_4800 replaced by ADD_11602

//ADD_4799 replaced by ADD_11602

//ADD_4798 replaced by ADD_11602

//ADD_4797 replaced by ADD_11602

//ADD_4796 replaced by ADD_11602

//ADD_4795 replaced by ADD_11602

//ADD_4794 replaced by ADD_11602

//ADD_4814 replaced by ADD_11601

//ADD_4813 replaced by ADD_11602

//ADD_4812 replaced by ADD_11602

//ADD_4811 replaced by ADD_11602

//ADD_4810 replaced by ADD_11602

//ADD_4809 replaced by ADD_11602

//ADD_4808 replaced by ADD_11602

//ADD_4807 replaced by ADD_11602

//ADD_4806 replaced by ADD_11602

//ADD_4822 replaced by ADD_11602

//ADD_4821 replaced by ADD_11602

//ADD_4820 replaced by ADD_11602

//ADD_4819 replaced by ADD_11602

//ADD_4818 replaced by ADD_11602

//ADD_4817 replaced by ADD_11602

//ADD_4816 replaced by ADD_11602

//ADD_4815 replaced by ADD_11602

//BADD_1435 replaced by BADD_1672

//BADD_1434 replaced by BADD_1671

//BADD_1433 replaced by BADD_1670

//ADD_4826 replaced by ADD_11602

//ADD_4825 replaced by ADD_11602

//ADD_4824 replaced by ADD_11602

//ADD_4823 replaced by ADD_11602

//KaratsubaCore_254 replaced by KaratsubaCore_467

//KaratsubaCore_253 replaced by KaratsubaCore_466

//KaratsubaCore_252 replaced by KaratsubaCore_465

//BADD_1439 replaced by BADD_1666

//BADD_1438 replaced by BADD_1668

//BADD_1437 replaced by BADD_1667

//BADD_1436 replaced by BADD_1666

//ADD_4830 replaced by ADD_8288

//ADD_4829 replaced by ADD_8288

//ADD_4828 replaced by ADD_8288

//ADD_4827 replaced by ADD_8288

//KaratsubaCore_257 replaced by KaratsubaCore_464

//KaratsubaCore_256 replaced by KaratsubaCore_463

//KaratsubaCore_255 replaced by KaratsubaCore_462

//BADD_1442 replaced by BADD_1672

//BADD_1441 replaced by BADD_1671

//BADD_1440 replaced by BADD_1670

//ADD_4834 replaced by ADD_11602

//ADD_4833 replaced by ADD_11602

//ADD_4832 replaced by ADD_11602

//ADD_4831 replaced by ADD_11602

//KaratsubaCore_260 replaced by KaratsubaCore_467

//KaratsubaCore_259 replaced by KaratsubaCore_466

//KaratsubaCore_258 replaced by KaratsubaCore_465

//ADD_4846 replaced by ADD_11602

//ADD_4845 replaced by ADD_11602

//ADD_4844 replaced by ADD_11602

//ADD_4843 replaced by ADD_11602

//ADD_4842 replaced by ADD_11602

//ADD_4841 replaced by ADD_11602

//ADD_4840 replaced by ADD_11602

//ADD_4839 replaced by ADD_11602

//ADD_4838 replaced by ADD_11602

//ADD_4837 replaced by ADD_11602

//ADD_4836 replaced by ADD_11602

//ADD_4835 replaced by ADD_11602

//ADD_4855 replaced by ADD_11601

//ADD_4854 replaced by ADD_11602

//ADD_4853 replaced by ADD_11602

//ADD_4852 replaced by ADD_11602

//ADD_4851 replaced by ADD_11602

//ADD_4850 replaced by ADD_11602

//ADD_4849 replaced by ADD_11602

//ADD_4848 replaced by ADD_11602

//ADD_4847 replaced by ADD_11602

//ADD_4863 replaced by ADD_11602

//ADD_4862 replaced by ADD_11602

//ADD_4861 replaced by ADD_11602

//ADD_4860 replaced by ADD_11602

//ADD_4859 replaced by ADD_11602

//ADD_4858 replaced by ADD_11602

//ADD_4857 replaced by ADD_11602

//ADD_4856 replaced by ADD_11602

//BADD_1445 replaced by BADD_1672

//BADD_1444 replaced by BADD_1671

//BADD_1443 replaced by BADD_1670

//ADD_4867 replaced by ADD_11602

//ADD_4866 replaced by ADD_11602

//ADD_4865 replaced by ADD_11602

//ADD_4864 replaced by ADD_11602

//KaratsubaCore_263 replaced by KaratsubaCore_467

//KaratsubaCore_262 replaced by KaratsubaCore_466

//KaratsubaCore_261 replaced by KaratsubaCore_465

//BADD_1449 replaced by BADD_1666

//BADD_1448 replaced by BADD_1668

//BADD_1447 replaced by BADD_1667

//BADD_1446 replaced by BADD_1666

//ADD_4871 replaced by ADD_8288

//ADD_4870 replaced by ADD_8288

//ADD_4869 replaced by ADD_8288

//ADD_4868 replaced by ADD_8288

//KaratsubaCore_266 replaced by KaratsubaCore_464

//KaratsubaCore_265 replaced by KaratsubaCore_463

//KaratsubaCore_264 replaced by KaratsubaCore_462

//BADD_1452 replaced by BADD_1672

//BADD_1451 replaced by BADD_1671

//BADD_1450 replaced by BADD_1670

//ADD_4875 replaced by ADD_11602

//ADD_4874 replaced by ADD_11602

//ADD_4873 replaced by ADD_11602

//ADD_4872 replaced by ADD_11602

//KaratsubaCore_269 replaced by KaratsubaCore_467

//KaratsubaCore_268 replaced by KaratsubaCore_466

//KaratsubaCore_267 replaced by KaratsubaCore_465

//ADD_4881 replaced by ADD_5761

//ADD_4880 replaced by ADD_5756

//ADD_4879 replaced by ADD_5756

//ADD_4878 replaced by ADD_5756

//ADD_4877 replaced by ADD_5756

//ADD_4876 replaced by ADD_5756

//ADD_4893 replaced by ADD_11602

//ADD_4892 replaced by ADD_11602

//ADD_4891 replaced by ADD_11602

//ADD_4890 replaced by ADD_11602

//ADD_4889 replaced by ADD_11602

//ADD_4888 replaced by ADD_11602

//ADD_4887 replaced by ADD_11602

//ADD_4886 replaced by ADD_11602

//ADD_4885 replaced by ADD_11602

//ADD_4884 replaced by ADD_11602

//ADD_4883 replaced by ADD_11602

//ADD_4882 replaced by ADD_11602

//ADD_4902 replaced by ADD_11601

//ADD_4901 replaced by ADD_11602

//ADD_4900 replaced by ADD_11602

//ADD_4899 replaced by ADD_11602

//ADD_4898 replaced by ADD_11602

//ADD_4897 replaced by ADD_11602

//ADD_4896 replaced by ADD_11602

//ADD_4895 replaced by ADD_11602

//ADD_4894 replaced by ADD_11602

//ADD_4910 replaced by ADD_11602

//ADD_4909 replaced by ADD_11602

//ADD_4908 replaced by ADD_11602

//ADD_4907 replaced by ADD_11602

//ADD_4906 replaced by ADD_11602

//ADD_4905 replaced by ADD_11602

//ADD_4904 replaced by ADD_11602

//ADD_4903 replaced by ADD_11602

//BADD_1455 replaced by BADD_1672

//BADD_1454 replaced by BADD_1671

//BADD_1453 replaced by BADD_1670

//ADD_4914 replaced by ADD_11602

//ADD_4913 replaced by ADD_11602

//ADD_4912 replaced by ADD_11602

//ADD_4911 replaced by ADD_11602

//KaratsubaCore_272 replaced by KaratsubaCore_467

//KaratsubaCore_271 replaced by KaratsubaCore_466

//KaratsubaCore_270 replaced by KaratsubaCore_465

//BADD_1459 replaced by BADD_1666

//BADD_1458 replaced by BADD_1668

//BADD_1457 replaced by BADD_1667

//BADD_1456 replaced by BADD_1666

//ADD_4918 replaced by ADD_8288

//ADD_4917 replaced by ADD_8288

//ADD_4916 replaced by ADD_8288

//ADD_4915 replaced by ADD_8288

//KaratsubaCore_275 replaced by KaratsubaCore_464

//KaratsubaCore_274 replaced by KaratsubaCore_463

//KaratsubaCore_273 replaced by KaratsubaCore_462

//BADD_1462 replaced by BADD_1672

//BADD_1461 replaced by BADD_1671

//BADD_1460 replaced by BADD_1670

//ADD_4922 replaced by ADD_11602

//ADD_4921 replaced by ADD_11602

//ADD_4920 replaced by ADD_11602

//ADD_4919 replaced by ADD_11602

//KaratsubaCore_278 replaced by KaratsubaCore_467

//KaratsubaCore_277 replaced by KaratsubaCore_466

//KaratsubaCore_276 replaced by KaratsubaCore_465

//ADD_4934 replaced by ADD_11602

//ADD_4933 replaced by ADD_11602

//ADD_4932 replaced by ADD_11602

//ADD_4931 replaced by ADD_11602

//ADD_4930 replaced by ADD_11602

//ADD_4929 replaced by ADD_11602

//ADD_4928 replaced by ADD_11602

//ADD_4927 replaced by ADD_11602

//ADD_4926 replaced by ADD_11602

//ADD_4925 replaced by ADD_11602

//ADD_4924 replaced by ADD_11602

//ADD_4923 replaced by ADD_11602

//ADD_4943 replaced by ADD_11601

//ADD_4942 replaced by ADD_11602

//ADD_4941 replaced by ADD_11602

//ADD_4940 replaced by ADD_11602

//ADD_4939 replaced by ADD_11602

//ADD_4938 replaced by ADD_11602

//ADD_4937 replaced by ADD_11602

//ADD_4936 replaced by ADD_11602

//ADD_4935 replaced by ADD_11602

//ADD_4951 replaced by ADD_11602

//ADD_4950 replaced by ADD_11602

//ADD_4949 replaced by ADD_11602

//ADD_4948 replaced by ADD_11602

//ADD_4947 replaced by ADD_11602

//ADD_4946 replaced by ADD_11602

//ADD_4945 replaced by ADD_11602

//ADD_4944 replaced by ADD_11602

//BADD_1465 replaced by BADD_1672

//BADD_1464 replaced by BADD_1671

//BADD_1463 replaced by BADD_1670

//ADD_4955 replaced by ADD_11602

//ADD_4954 replaced by ADD_11602

//ADD_4953 replaced by ADD_11602

//ADD_4952 replaced by ADD_11602

//KaratsubaCore_281 replaced by KaratsubaCore_467

//KaratsubaCore_280 replaced by KaratsubaCore_466

//KaratsubaCore_279 replaced by KaratsubaCore_465

//BADD_1469 replaced by BADD_1666

//BADD_1468 replaced by BADD_1668

//BADD_1467 replaced by BADD_1667

//BADD_1466 replaced by BADD_1666

//ADD_4959 replaced by ADD_8288

//ADD_4958 replaced by ADD_8288

//ADD_4957 replaced by ADD_8288

//ADD_4956 replaced by ADD_8288

//KaratsubaCore_284 replaced by KaratsubaCore_464

//KaratsubaCore_283 replaced by KaratsubaCore_463

//KaratsubaCore_282 replaced by KaratsubaCore_462

//BADD_1472 replaced by BADD_1672

//BADD_1471 replaced by BADD_1671

//BADD_1470 replaced by BADD_1670

//ADD_4963 replaced by ADD_11602

//ADD_4962 replaced by ADD_11602

//ADD_4961 replaced by ADD_11602

//ADD_4960 replaced by ADD_11602

//KaratsubaCore_287 replaced by KaratsubaCore_467

//KaratsubaCore_286 replaced by KaratsubaCore_466

//KaratsubaCore_285 replaced by KaratsubaCore_465

//ADD_4969 replaced by ADD_5761

//ADD_4968 replaced by ADD_5756

//ADD_4967 replaced by ADD_5756

//ADD_4966 replaced by ADD_5756

//ADD_4965 replaced by ADD_5756

//ADD_4964 replaced by ADD_5756

//ADD_4981 replaced by ADD_11602

//ADD_4980 replaced by ADD_11602

//ADD_4979 replaced by ADD_11602

//ADD_4978 replaced by ADD_11602

//ADD_4977 replaced by ADD_11602

//ADD_4976 replaced by ADD_11602

//ADD_4975 replaced by ADD_11602

//ADD_4974 replaced by ADD_11602

//ADD_4973 replaced by ADD_11602

//ADD_4972 replaced by ADD_11602

//ADD_4971 replaced by ADD_11602

//ADD_4970 replaced by ADD_11602

//ADD_4990 replaced by ADD_11601

//ADD_4989 replaced by ADD_11602

//ADD_4988 replaced by ADD_11602

//ADD_4987 replaced by ADD_11602

//ADD_4986 replaced by ADD_11602

//ADD_4985 replaced by ADD_11602

//ADD_4984 replaced by ADD_11602

//ADD_4983 replaced by ADD_11602

//ADD_4982 replaced by ADD_11602

//ADD_4998 replaced by ADD_11602

//ADD_4997 replaced by ADD_11602

//ADD_4996 replaced by ADD_11602

//ADD_4995 replaced by ADD_11602

//ADD_4994 replaced by ADD_11602

//ADD_4993 replaced by ADD_11602

//ADD_4992 replaced by ADD_11602

//ADD_4991 replaced by ADD_11602

//BADD_1475 replaced by BADD_1672

//BADD_1474 replaced by BADD_1671

//BADD_1473 replaced by BADD_1670

//ADD_5002 replaced by ADD_11602

//ADD_5001 replaced by ADD_11602

//ADD_5000 replaced by ADD_11602

//ADD_4999 replaced by ADD_11602

//KaratsubaCore_290 replaced by KaratsubaCore_467

//KaratsubaCore_289 replaced by KaratsubaCore_466

//KaratsubaCore_288 replaced by KaratsubaCore_465

//BADD_1479 replaced by BADD_1666

//BADD_1478 replaced by BADD_1668

//BADD_1477 replaced by BADD_1667

//BADD_1476 replaced by BADD_1666

//ADD_5006 replaced by ADD_8288

//ADD_5005 replaced by ADD_8288

//ADD_5004 replaced by ADD_8288

//ADD_5003 replaced by ADD_8288

//KaratsubaCore_293 replaced by KaratsubaCore_464

//KaratsubaCore_292 replaced by KaratsubaCore_463

//KaratsubaCore_291 replaced by KaratsubaCore_462

//BADD_1482 replaced by BADD_1672

//BADD_1481 replaced by BADD_1671

//BADD_1480 replaced by BADD_1670

//ADD_5010 replaced by ADD_11602

//ADD_5009 replaced by ADD_11602

//ADD_5008 replaced by ADD_11602

//ADD_5007 replaced by ADD_11602

//KaratsubaCore_296 replaced by KaratsubaCore_467

//KaratsubaCore_295 replaced by KaratsubaCore_466

//KaratsubaCore_294 replaced by KaratsubaCore_465

//ADD_5022 replaced by ADD_11602

//ADD_5021 replaced by ADD_11602

//ADD_5020 replaced by ADD_11602

//ADD_5019 replaced by ADD_11602

//ADD_5018 replaced by ADD_11602

//ADD_5017 replaced by ADD_11602

//ADD_5016 replaced by ADD_11602

//ADD_5015 replaced by ADD_11602

//ADD_5014 replaced by ADD_11602

//ADD_5013 replaced by ADD_11602

//ADD_5012 replaced by ADD_11602

//ADD_5011 replaced by ADD_11602

//ADD_5031 replaced by ADD_11601

//ADD_5030 replaced by ADD_11602

//ADD_5029 replaced by ADD_11602

//ADD_5028 replaced by ADD_11602

//ADD_5027 replaced by ADD_11602

//ADD_5026 replaced by ADD_11602

//ADD_5025 replaced by ADD_11602

//ADD_5024 replaced by ADD_11602

//ADD_5023 replaced by ADD_11602

//ADD_5039 replaced by ADD_11602

//ADD_5038 replaced by ADD_11602

//ADD_5037 replaced by ADD_11602

//ADD_5036 replaced by ADD_11602

//ADD_5035 replaced by ADD_11602

//ADD_5034 replaced by ADD_11602

//ADD_5033 replaced by ADD_11602

//ADD_5032 replaced by ADD_11602

//BADD_1485 replaced by BADD_1672

//BADD_1484 replaced by BADD_1671

//BADD_1483 replaced by BADD_1670

//ADD_5043 replaced by ADD_11602

//ADD_5042 replaced by ADD_11602

//ADD_5041 replaced by ADD_11602

//ADD_5040 replaced by ADD_11602

//KaratsubaCore_299 replaced by KaratsubaCore_467

//KaratsubaCore_298 replaced by KaratsubaCore_466

//KaratsubaCore_297 replaced by KaratsubaCore_465

//BADD_1489 replaced by BADD_1666

//BADD_1488 replaced by BADD_1668

//BADD_1487 replaced by BADD_1667

//BADD_1486 replaced by BADD_1666

//ADD_5047 replaced by ADD_8288

//ADD_5046 replaced by ADD_8288

//ADD_5045 replaced by ADD_8288

//ADD_5044 replaced by ADD_8288

//KaratsubaCore_302 replaced by KaratsubaCore_464

//KaratsubaCore_301 replaced by KaratsubaCore_463

//KaratsubaCore_300 replaced by KaratsubaCore_462

//BADD_1492 replaced by BADD_1672

//BADD_1491 replaced by BADD_1671

//BADD_1490 replaced by BADD_1670

//ADD_5051 replaced by ADD_11602

//ADD_5050 replaced by ADD_11602

//ADD_5049 replaced by ADD_11602

//ADD_5048 replaced by ADD_11602

//KaratsubaCore_305 replaced by KaratsubaCore_467

//KaratsubaCore_304 replaced by KaratsubaCore_466

//KaratsubaCore_303 replaced by KaratsubaCore_465

//ADD_5057 replaced by ADD_5761

//ADD_5056 replaced by ADD_5756

//ADD_5055 replaced by ADD_5756

//ADD_5054 replaced by ADD_5756

//ADD_5053 replaced by ADD_5756

//ADD_5052 replaced by ADD_5756

//ADD_5069 replaced by ADD_11602

//ADD_5068 replaced by ADD_11602

//ADD_5067 replaced by ADD_11602

//ADD_5066 replaced by ADD_11602

//ADD_5065 replaced by ADD_11602

//ADD_5064 replaced by ADD_11602

//ADD_5063 replaced by ADD_11602

//ADD_5062 replaced by ADD_11602

//ADD_5061 replaced by ADD_11602

//ADD_5060 replaced by ADD_11602

//ADD_5059 replaced by ADD_11602

//ADD_5058 replaced by ADD_11602

//ADD_5078 replaced by ADD_11601

//ADD_5077 replaced by ADD_11602

//ADD_5076 replaced by ADD_11602

//ADD_5075 replaced by ADD_11602

//ADD_5074 replaced by ADD_11602

//ADD_5073 replaced by ADD_11602

//ADD_5072 replaced by ADD_11602

//ADD_5071 replaced by ADD_11602

//ADD_5070 replaced by ADD_11602

//ADD_5086 replaced by ADD_11602

//ADD_5085 replaced by ADD_11602

//ADD_5084 replaced by ADD_11602

//ADD_5083 replaced by ADD_11602

//ADD_5082 replaced by ADD_11602

//ADD_5081 replaced by ADD_11602

//ADD_5080 replaced by ADD_11602

//ADD_5079 replaced by ADD_11602

//BADD_1495 replaced by BADD_1672

//BADD_1494 replaced by BADD_1671

//BADD_1493 replaced by BADD_1670

//ADD_5090 replaced by ADD_11602

//ADD_5089 replaced by ADD_11602

//ADD_5088 replaced by ADD_11602

//ADD_5087 replaced by ADD_11602

//KaratsubaCore_308 replaced by KaratsubaCore_467

//KaratsubaCore_307 replaced by KaratsubaCore_466

//KaratsubaCore_306 replaced by KaratsubaCore_465

//BADD_1499 replaced by BADD_1666

//BADD_1498 replaced by BADD_1668

//BADD_1497 replaced by BADD_1667

//BADD_1496 replaced by BADD_1666

//ADD_5094 replaced by ADD_8288

//ADD_5093 replaced by ADD_8288

//ADD_5092 replaced by ADD_8288

//ADD_5091 replaced by ADD_8288

//KaratsubaCore_311 replaced by KaratsubaCore_464

//KaratsubaCore_310 replaced by KaratsubaCore_463

//KaratsubaCore_309 replaced by KaratsubaCore_462

//BADD_1502 replaced by BADD_1672

//BADD_1501 replaced by BADD_1671

//BADD_1500 replaced by BADD_1670

//ADD_5098 replaced by ADD_11602

//ADD_5097 replaced by ADD_11602

//ADD_5096 replaced by ADD_11602

//ADD_5095 replaced by ADD_11602

//KaratsubaCore_314 replaced by KaratsubaCore_467

//KaratsubaCore_313 replaced by KaratsubaCore_466

//KaratsubaCore_312 replaced by KaratsubaCore_465

//ADD_5110 replaced by ADD_11602

//ADD_5109 replaced by ADD_11602

//ADD_5108 replaced by ADD_11602

//ADD_5107 replaced by ADD_11602

//ADD_5106 replaced by ADD_11602

//ADD_5105 replaced by ADD_11602

//ADD_5104 replaced by ADD_11602

//ADD_5103 replaced by ADD_11602

//ADD_5102 replaced by ADD_11602

//ADD_5101 replaced by ADD_11602

//ADD_5100 replaced by ADD_11602

//ADD_5099 replaced by ADD_11602

//ADD_5119 replaced by ADD_11601

//ADD_5118 replaced by ADD_11602

//ADD_5117 replaced by ADD_11602

//ADD_5116 replaced by ADD_11602

//ADD_5115 replaced by ADD_11602

//ADD_5114 replaced by ADD_11602

//ADD_5113 replaced by ADD_11602

//ADD_5112 replaced by ADD_11602

//ADD_5111 replaced by ADD_11602

//ADD_5127 replaced by ADD_11602

//ADD_5126 replaced by ADD_11602

//ADD_5125 replaced by ADD_11602

//ADD_5124 replaced by ADD_11602

//ADD_5123 replaced by ADD_11602

//ADD_5122 replaced by ADD_11602

//ADD_5121 replaced by ADD_11602

//ADD_5120 replaced by ADD_11602

//BADD_1505 replaced by BADD_1672

//BADD_1504 replaced by BADD_1671

//BADD_1503 replaced by BADD_1670

//ADD_5131 replaced by ADD_11602

//ADD_5130 replaced by ADD_11602

//ADD_5129 replaced by ADD_11602

//ADD_5128 replaced by ADD_11602

//KaratsubaCore_317 replaced by KaratsubaCore_467

//KaratsubaCore_316 replaced by KaratsubaCore_466

//KaratsubaCore_315 replaced by KaratsubaCore_465

//BADD_1509 replaced by BADD_1666

//BADD_1508 replaced by BADD_1668

//BADD_1507 replaced by BADD_1667

//BADD_1506 replaced by BADD_1666

//ADD_5135 replaced by ADD_8288

//ADD_5134 replaced by ADD_8288

//ADD_5133 replaced by ADD_8288

//ADD_5132 replaced by ADD_8288

//KaratsubaCore_320 replaced by KaratsubaCore_464

//KaratsubaCore_319 replaced by KaratsubaCore_463

//KaratsubaCore_318 replaced by KaratsubaCore_462

//BADD_1512 replaced by BADD_1672

//BADD_1511 replaced by BADD_1671

//BADD_1510 replaced by BADD_1670

//ADD_5139 replaced by ADD_11602

//ADD_5138 replaced by ADD_11602

//ADD_5137 replaced by ADD_11602

//ADD_5136 replaced by ADD_11602

//KaratsubaCore_323 replaced by KaratsubaCore_467

//KaratsubaCore_322 replaced by KaratsubaCore_466

//KaratsubaCore_321 replaced by KaratsubaCore_465

//ADD_5145 replaced by ADD_5761

//ADD_5144 replaced by ADD_5756

//ADD_5143 replaced by ADD_5756

//ADD_5142 replaced by ADD_5756

//ADD_5141 replaced by ADD_5756

//ADD_5140 replaced by ADD_5756

//ADD_5157 replaced by ADD_11602

//ADD_5156 replaced by ADD_11602

//ADD_5155 replaced by ADD_11602

//ADD_5154 replaced by ADD_11602

//ADD_5153 replaced by ADD_11602

//ADD_5152 replaced by ADD_11602

//ADD_5151 replaced by ADD_11602

//ADD_5150 replaced by ADD_11602

//ADD_5149 replaced by ADD_11602

//ADD_5148 replaced by ADD_11602

//ADD_5147 replaced by ADD_11602

//ADD_5146 replaced by ADD_11602

//ADD_5166 replaced by ADD_11601

//ADD_5165 replaced by ADD_11602

//ADD_5164 replaced by ADD_11602

//ADD_5163 replaced by ADD_11602

//ADD_5162 replaced by ADD_11602

//ADD_5161 replaced by ADD_11602

//ADD_5160 replaced by ADD_11602

//ADD_5159 replaced by ADD_11602

//ADD_5158 replaced by ADD_11602

//ADD_5174 replaced by ADD_11602

//ADD_5173 replaced by ADD_11602

//ADD_5172 replaced by ADD_11602

//ADD_5171 replaced by ADD_11602

//ADD_5170 replaced by ADD_11602

//ADD_5169 replaced by ADD_11602

//ADD_5168 replaced by ADD_11602

//ADD_5167 replaced by ADD_11602

//BADD_1515 replaced by BADD_1672

//BADD_1514 replaced by BADD_1671

//BADD_1513 replaced by BADD_1670

//ADD_5178 replaced by ADD_11602

//ADD_5177 replaced by ADD_11602

//ADD_5176 replaced by ADD_11602

//ADD_5175 replaced by ADD_11602

//KaratsubaCore_326 replaced by KaratsubaCore_467

//KaratsubaCore_325 replaced by KaratsubaCore_466

//KaratsubaCore_324 replaced by KaratsubaCore_465

//BADD_1519 replaced by BADD_1666

//BADD_1518 replaced by BADD_1668

//BADD_1517 replaced by BADD_1667

//BADD_1516 replaced by BADD_1666

//ADD_5182 replaced by ADD_8288

//ADD_5181 replaced by ADD_8288

//ADD_5180 replaced by ADD_8288

//ADD_5179 replaced by ADD_8288

//KaratsubaCore_329 replaced by KaratsubaCore_464

//KaratsubaCore_328 replaced by KaratsubaCore_463

//KaratsubaCore_327 replaced by KaratsubaCore_462

//BADD_1522 replaced by BADD_1672

//BADD_1521 replaced by BADD_1671

//BADD_1520 replaced by BADD_1670

//ADD_5186 replaced by ADD_11602

//ADD_5185 replaced by ADD_11602

//ADD_5184 replaced by ADD_11602

//ADD_5183 replaced by ADD_11602

//KaratsubaCore_332 replaced by KaratsubaCore_467

//KaratsubaCore_331 replaced by KaratsubaCore_466

//KaratsubaCore_330 replaced by KaratsubaCore_465

//ADD_5198 replaced by ADD_11602

//ADD_5197 replaced by ADD_11602

//ADD_5196 replaced by ADD_11602

//ADD_5195 replaced by ADD_11602

//ADD_5194 replaced by ADD_11602

//ADD_5193 replaced by ADD_11602

//ADD_5192 replaced by ADD_11602

//ADD_5191 replaced by ADD_11602

//ADD_5190 replaced by ADD_11602

//ADD_5189 replaced by ADD_11602

//ADD_5188 replaced by ADD_11602

//ADD_5187 replaced by ADD_11602

//ADD_5207 replaced by ADD_11601

//ADD_5206 replaced by ADD_11602

//ADD_5205 replaced by ADD_11602

//ADD_5204 replaced by ADD_11602

//ADD_5203 replaced by ADD_11602

//ADD_5202 replaced by ADD_11602

//ADD_5201 replaced by ADD_11602

//ADD_5200 replaced by ADD_11602

//ADD_5199 replaced by ADD_11602

//ADD_5215 replaced by ADD_11602

//ADD_5214 replaced by ADD_11602

//ADD_5213 replaced by ADD_11602

//ADD_5212 replaced by ADD_11602

//ADD_5211 replaced by ADD_11602

//ADD_5210 replaced by ADD_11602

//ADD_5209 replaced by ADD_11602

//ADD_5208 replaced by ADD_11602

//BADD_1525 replaced by BADD_1672

//BADD_1524 replaced by BADD_1671

//BADD_1523 replaced by BADD_1670

//ADD_5219 replaced by ADD_11602

//ADD_5218 replaced by ADD_11602

//ADD_5217 replaced by ADD_11602

//ADD_5216 replaced by ADD_11602

//KaratsubaCore_335 replaced by KaratsubaCore_467

//KaratsubaCore_334 replaced by KaratsubaCore_466

//KaratsubaCore_333 replaced by KaratsubaCore_465

//BADD_1529 replaced by BADD_1666

//BADD_1528 replaced by BADD_1668

//BADD_1527 replaced by BADD_1667

//BADD_1526 replaced by BADD_1666

//ADD_5223 replaced by ADD_8288

//ADD_5222 replaced by ADD_8288

//ADD_5221 replaced by ADD_8288

//ADD_5220 replaced by ADD_8288

//KaratsubaCore_338 replaced by KaratsubaCore_464

//KaratsubaCore_337 replaced by KaratsubaCore_463

//KaratsubaCore_336 replaced by KaratsubaCore_462

//BADD_1532 replaced by BADD_1672

//BADD_1531 replaced by BADD_1671

//BADD_1530 replaced by BADD_1670

//ADD_5227 replaced by ADD_11602

//ADD_5226 replaced by ADD_11602

//ADD_5225 replaced by ADD_11602

//ADD_5224 replaced by ADD_11602

//KaratsubaCore_341 replaced by KaratsubaCore_467

//KaratsubaCore_340 replaced by KaratsubaCore_466

//KaratsubaCore_339 replaced by KaratsubaCore_465

//ADD_5233 replaced by ADD_5761

//ADD_5232 replaced by ADD_5756

//ADD_5231 replaced by ADD_5756

//ADD_5230 replaced by ADD_5756

//ADD_5229 replaced by ADD_5756

//ADD_5228 replaced by ADD_5756

//ADD_5245 replaced by ADD_11602

//ADD_5244 replaced by ADD_11602

//ADD_5243 replaced by ADD_11602

//ADD_5242 replaced by ADD_11602

//ADD_5241 replaced by ADD_11602

//ADD_5240 replaced by ADD_11602

//ADD_5239 replaced by ADD_11602

//ADD_5238 replaced by ADD_11602

//ADD_5237 replaced by ADD_11602

//ADD_5236 replaced by ADD_11602

//ADD_5235 replaced by ADD_11602

//ADD_5234 replaced by ADD_11602

//ADD_5254 replaced by ADD_11601

//ADD_5253 replaced by ADD_11602

//ADD_5252 replaced by ADD_11602

//ADD_5251 replaced by ADD_11602

//ADD_5250 replaced by ADD_11602

//ADD_5249 replaced by ADD_11602

//ADD_5248 replaced by ADD_11602

//ADD_5247 replaced by ADD_11602

//ADD_5246 replaced by ADD_11602

//ADD_5262 replaced by ADD_11602

//ADD_5261 replaced by ADD_11602

//ADD_5260 replaced by ADD_11602

//ADD_5259 replaced by ADD_11602

//ADD_5258 replaced by ADD_11602

//ADD_5257 replaced by ADD_11602

//ADD_5256 replaced by ADD_11602

//ADD_5255 replaced by ADD_11602

//BADD_1535 replaced by BADD_1672

//BADD_1534 replaced by BADD_1671

//BADD_1533 replaced by BADD_1670

//ADD_5266 replaced by ADD_11602

//ADD_5265 replaced by ADD_11602

//ADD_5264 replaced by ADD_11602

//ADD_5263 replaced by ADD_11602

//KaratsubaCore_344 replaced by KaratsubaCore_467

//KaratsubaCore_343 replaced by KaratsubaCore_466

//KaratsubaCore_342 replaced by KaratsubaCore_465

//BADD_1539 replaced by BADD_1666

//BADD_1538 replaced by BADD_1668

//BADD_1537 replaced by BADD_1667

//BADD_1536 replaced by BADD_1666

//ADD_5270 replaced by ADD_8288

//ADD_5269 replaced by ADD_8288

//ADD_5268 replaced by ADD_8288

//ADD_5267 replaced by ADD_8288

//KaratsubaCore_347 replaced by KaratsubaCore_464

//KaratsubaCore_346 replaced by KaratsubaCore_463

//KaratsubaCore_345 replaced by KaratsubaCore_462

//BADD_1542 replaced by BADD_1672

//BADD_1541 replaced by BADD_1671

//BADD_1540 replaced by BADD_1670

//ADD_5274 replaced by ADD_11602

//ADD_5273 replaced by ADD_11602

//ADD_5272 replaced by ADD_11602

//ADD_5271 replaced by ADD_11602

//KaratsubaCore_350 replaced by KaratsubaCore_467

//KaratsubaCore_349 replaced by KaratsubaCore_466

//KaratsubaCore_348 replaced by KaratsubaCore_465

//ADD_5286 replaced by ADD_11602

//ADD_5285 replaced by ADD_11602

//ADD_5284 replaced by ADD_11602

//ADD_5283 replaced by ADD_11602

//ADD_5282 replaced by ADD_11602

//ADD_5281 replaced by ADD_11602

//ADD_5280 replaced by ADD_11602

//ADD_5279 replaced by ADD_11602

//ADD_5278 replaced by ADD_11602

//ADD_5277 replaced by ADD_11602

//ADD_5276 replaced by ADD_11602

//ADD_5275 replaced by ADD_11602

//ADD_5295 replaced by ADD_11601

//ADD_5294 replaced by ADD_11602

//ADD_5293 replaced by ADD_11602

//ADD_5292 replaced by ADD_11602

//ADD_5291 replaced by ADD_11602

//ADD_5290 replaced by ADD_11602

//ADD_5289 replaced by ADD_11602

//ADD_5288 replaced by ADD_11602

//ADD_5287 replaced by ADD_11602

//ADD_5303 replaced by ADD_11602

//ADD_5302 replaced by ADD_11602

//ADD_5301 replaced by ADD_11602

//ADD_5300 replaced by ADD_11602

//ADD_5299 replaced by ADD_11602

//ADD_5298 replaced by ADD_11602

//ADD_5297 replaced by ADD_11602

//ADD_5296 replaced by ADD_11602

//BADD_1545 replaced by BADD_1672

//BADD_1544 replaced by BADD_1671

//BADD_1543 replaced by BADD_1670

//ADD_5307 replaced by ADD_11602

//ADD_5306 replaced by ADD_11602

//ADD_5305 replaced by ADD_11602

//ADD_5304 replaced by ADD_11602

//KaratsubaCore_353 replaced by KaratsubaCore_467

//KaratsubaCore_352 replaced by KaratsubaCore_466

//KaratsubaCore_351 replaced by KaratsubaCore_465

//BADD_1549 replaced by BADD_1666

//BADD_1548 replaced by BADD_1668

//BADD_1547 replaced by BADD_1667

//BADD_1546 replaced by BADD_1666

//ADD_5311 replaced by ADD_8288

//ADD_5310 replaced by ADD_8288

//ADD_5309 replaced by ADD_8288

//ADD_5308 replaced by ADD_8288

//KaratsubaCore_356 replaced by KaratsubaCore_464

//KaratsubaCore_355 replaced by KaratsubaCore_463

//KaratsubaCore_354 replaced by KaratsubaCore_462

//BADD_1552 replaced by BADD_1672

//BADD_1551 replaced by BADD_1671

//BADD_1550 replaced by BADD_1670

//ADD_5315 replaced by ADD_11602

//ADD_5314 replaced by ADD_11602

//ADD_5313 replaced by ADD_11602

//ADD_5312 replaced by ADD_11602

//KaratsubaCore_359 replaced by KaratsubaCore_467

//KaratsubaCore_358 replaced by KaratsubaCore_466

//KaratsubaCore_357 replaced by KaratsubaCore_465

//ADD_5321 replaced by ADD_5761

//ADD_5320 replaced by ADD_5756

//ADD_5319 replaced by ADD_5756

//ADD_5318 replaced by ADD_5756

//ADD_5317 replaced by ADD_5756

//ADD_5316 replaced by ADD_5756

//ADD_5333 replaced by ADD_11602

//ADD_5332 replaced by ADD_11602

//ADD_5331 replaced by ADD_11602

//ADD_5330 replaced by ADD_11602

//ADD_5329 replaced by ADD_11602

//ADD_5328 replaced by ADD_11602

//ADD_5327 replaced by ADD_11602

//ADD_5326 replaced by ADD_11602

//ADD_5325 replaced by ADD_11602

//ADD_5324 replaced by ADD_11602

//ADD_5323 replaced by ADD_11602

//ADD_5322 replaced by ADD_11602

//ADD_5342 replaced by ADD_11601

//ADD_5341 replaced by ADD_11602

//ADD_5340 replaced by ADD_11602

//ADD_5339 replaced by ADD_11602

//ADD_5338 replaced by ADD_11602

//ADD_5337 replaced by ADD_11602

//ADD_5336 replaced by ADD_11602

//ADD_5335 replaced by ADD_11602

//ADD_5334 replaced by ADD_11602

//ADD_5350 replaced by ADD_11602

//ADD_5349 replaced by ADD_11602

//ADD_5348 replaced by ADD_11602

//ADD_5347 replaced by ADD_11602

//ADD_5346 replaced by ADD_11602

//ADD_5345 replaced by ADD_11602

//ADD_5344 replaced by ADD_11602

//ADD_5343 replaced by ADD_11602

//BADD_1555 replaced by BADD_1672

//BADD_1554 replaced by BADD_1671

//BADD_1553 replaced by BADD_1670

//ADD_5354 replaced by ADD_11602

//ADD_5353 replaced by ADD_11602

//ADD_5352 replaced by ADD_11602

//ADD_5351 replaced by ADD_11602

//KaratsubaCore_362 replaced by KaratsubaCore_467

//KaratsubaCore_361 replaced by KaratsubaCore_466

//KaratsubaCore_360 replaced by KaratsubaCore_465

//BADD_1559 replaced by BADD_1666

//BADD_1558 replaced by BADD_1668

//BADD_1557 replaced by BADD_1667

//BADD_1556 replaced by BADD_1666

//ADD_5358 replaced by ADD_8288

//ADD_5357 replaced by ADD_8288

//ADD_5356 replaced by ADD_8288

//ADD_5355 replaced by ADD_8288

//KaratsubaCore_365 replaced by KaratsubaCore_464

//KaratsubaCore_364 replaced by KaratsubaCore_463

//KaratsubaCore_363 replaced by KaratsubaCore_462

//BADD_1562 replaced by BADD_1672

//BADD_1561 replaced by BADD_1671

//BADD_1560 replaced by BADD_1670

//ADD_5362 replaced by ADD_11602

//ADD_5361 replaced by ADD_11602

//ADD_5360 replaced by ADD_11602

//ADD_5359 replaced by ADD_11602

//KaratsubaCore_368 replaced by KaratsubaCore_467

//KaratsubaCore_367 replaced by KaratsubaCore_466

//KaratsubaCore_366 replaced by KaratsubaCore_465

//ADD_5374 replaced by ADD_11602

//ADD_5373 replaced by ADD_11602

//ADD_5372 replaced by ADD_11602

//ADD_5371 replaced by ADD_11602

//ADD_5370 replaced by ADD_11602

//ADD_5369 replaced by ADD_11602

//ADD_5368 replaced by ADD_11602

//ADD_5367 replaced by ADD_11602

//ADD_5366 replaced by ADD_11602

//ADD_5365 replaced by ADD_11602

//ADD_5364 replaced by ADD_11602

//ADD_5363 replaced by ADD_11602

//ADD_5383 replaced by ADD_11601

//ADD_5382 replaced by ADD_11602

//ADD_5381 replaced by ADD_11602

//ADD_5380 replaced by ADD_11602

//ADD_5379 replaced by ADD_11602

//ADD_5378 replaced by ADD_11602

//ADD_5377 replaced by ADD_11602

//ADD_5376 replaced by ADD_11602

//ADD_5375 replaced by ADD_11602

//ADD_5391 replaced by ADD_11602

//ADD_5390 replaced by ADD_11602

//ADD_5389 replaced by ADD_11602

//ADD_5388 replaced by ADD_11602

//ADD_5387 replaced by ADD_11602

//ADD_5386 replaced by ADD_11602

//ADD_5385 replaced by ADD_11602

//ADD_5384 replaced by ADD_11602

//BADD_1565 replaced by BADD_1672

//BADD_1564 replaced by BADD_1671

//BADD_1563 replaced by BADD_1670

//ADD_5395 replaced by ADD_11602

//ADD_5394 replaced by ADD_11602

//ADD_5393 replaced by ADD_11602

//ADD_5392 replaced by ADD_11602

//KaratsubaCore_371 replaced by KaratsubaCore_467

//KaratsubaCore_370 replaced by KaratsubaCore_466

//KaratsubaCore_369 replaced by KaratsubaCore_465

//BADD_1569 replaced by BADD_1666

//BADD_1568 replaced by BADD_1668

//BADD_1567 replaced by BADD_1667

//BADD_1566 replaced by BADD_1666

//ADD_5399 replaced by ADD_8288

//ADD_5398 replaced by ADD_8288

//ADD_5397 replaced by ADD_8288

//ADD_5396 replaced by ADD_8288

//KaratsubaCore_374 replaced by KaratsubaCore_464

//KaratsubaCore_373 replaced by KaratsubaCore_463

//KaratsubaCore_372 replaced by KaratsubaCore_462

//BADD_1572 replaced by BADD_1672

//BADD_1571 replaced by BADD_1671

//BADD_1570 replaced by BADD_1670

//ADD_5403 replaced by ADD_11602

//ADD_5402 replaced by ADD_11602

//ADD_5401 replaced by ADD_11602

//ADD_5400 replaced by ADD_11602

//KaratsubaCore_377 replaced by KaratsubaCore_467

//KaratsubaCore_376 replaced by KaratsubaCore_466

//KaratsubaCore_375 replaced by KaratsubaCore_465

//ADD_5409 replaced by ADD_5761

//ADD_5408 replaced by ADD_5756

//ADD_5407 replaced by ADD_5756

//ADD_5406 replaced by ADD_5756

//ADD_5405 replaced by ADD_5756

//ADD_5404 replaced by ADD_5756

//ADD_5421 replaced by ADD_11602

//ADD_5420 replaced by ADD_11602

//ADD_5419 replaced by ADD_11602

//ADD_5418 replaced by ADD_11602

//ADD_5417 replaced by ADD_11602

//ADD_5416 replaced by ADD_11602

//ADD_5415 replaced by ADD_11602

//ADD_5414 replaced by ADD_11602

//ADD_5413 replaced by ADD_11602

//ADD_5412 replaced by ADD_11602

//ADD_5411 replaced by ADD_11602

//ADD_5410 replaced by ADD_11602

//ADD_5430 replaced by ADD_11601

//ADD_5429 replaced by ADD_11602

//ADD_5428 replaced by ADD_11602

//ADD_5427 replaced by ADD_11602

//ADD_5426 replaced by ADD_11602

//ADD_5425 replaced by ADD_11602

//ADD_5424 replaced by ADD_11602

//ADD_5423 replaced by ADD_11602

//ADD_5422 replaced by ADD_11602

//ADD_5438 replaced by ADD_11602

//ADD_5437 replaced by ADD_11602

//ADD_5436 replaced by ADD_11602

//ADD_5435 replaced by ADD_11602

//ADD_5434 replaced by ADD_11602

//ADD_5433 replaced by ADD_11602

//ADD_5432 replaced by ADD_11602

//ADD_5431 replaced by ADD_11602

//BADD_1575 replaced by BADD_1672

//BADD_1574 replaced by BADD_1671

//BADD_1573 replaced by BADD_1670

//ADD_5442 replaced by ADD_11602

//ADD_5441 replaced by ADD_11602

//ADD_5440 replaced by ADD_11602

//ADD_5439 replaced by ADD_11602

//KaratsubaCore_380 replaced by KaratsubaCore_467

//KaratsubaCore_379 replaced by KaratsubaCore_466

//KaratsubaCore_378 replaced by KaratsubaCore_465

//BADD_1579 replaced by BADD_1666

//BADD_1578 replaced by BADD_1668

//BADD_1577 replaced by BADD_1667

//BADD_1576 replaced by BADD_1666

//ADD_5446 replaced by ADD_8288

//ADD_5445 replaced by ADD_8288

//ADD_5444 replaced by ADD_8288

//ADD_5443 replaced by ADD_8288

//KaratsubaCore_383 replaced by KaratsubaCore_464

//KaratsubaCore_382 replaced by KaratsubaCore_463

//KaratsubaCore_381 replaced by KaratsubaCore_462

//BADD_1582 replaced by BADD_1672

//BADD_1581 replaced by BADD_1671

//BADD_1580 replaced by BADD_1670

//ADD_5450 replaced by ADD_11602

//ADD_5449 replaced by ADD_11602

//ADD_5448 replaced by ADD_11602

//ADD_5447 replaced by ADD_11602

//KaratsubaCore_386 replaced by KaratsubaCore_467

//KaratsubaCore_385 replaced by KaratsubaCore_466

//KaratsubaCore_384 replaced by KaratsubaCore_465

//ADD_5462 replaced by ADD_11602

//ADD_5461 replaced by ADD_11602

//ADD_5460 replaced by ADD_11602

//ADD_5459 replaced by ADD_11602

//ADD_5458 replaced by ADD_11602

//ADD_5457 replaced by ADD_11602

//ADD_5456 replaced by ADD_11602

//ADD_5455 replaced by ADD_11602

//ADD_5454 replaced by ADD_11602

//ADD_5453 replaced by ADD_11602

//ADD_5452 replaced by ADD_11602

//ADD_5451 replaced by ADD_11602

//ADD_5471 replaced by ADD_11601

//ADD_5470 replaced by ADD_11602

//ADD_5469 replaced by ADD_11602

//ADD_5468 replaced by ADD_11602

//ADD_5467 replaced by ADD_11602

//ADD_5466 replaced by ADD_11602

//ADD_5465 replaced by ADD_11602

//ADD_5464 replaced by ADD_11602

//ADD_5463 replaced by ADD_11602

//ADD_5479 replaced by ADD_11602

//ADD_5478 replaced by ADD_11602

//ADD_5477 replaced by ADD_11602

//ADD_5476 replaced by ADD_11602

//ADD_5475 replaced by ADD_11602

//ADD_5474 replaced by ADD_11602

//ADD_5473 replaced by ADD_11602

//ADD_5472 replaced by ADD_11602

//BADD_1585 replaced by BADD_1672

//BADD_1584 replaced by BADD_1671

//BADD_1583 replaced by BADD_1670

//ADD_5483 replaced by ADD_11602

//ADD_5482 replaced by ADD_11602

//ADD_5481 replaced by ADD_11602

//ADD_5480 replaced by ADD_11602

//KaratsubaCore_389 replaced by KaratsubaCore_467

//KaratsubaCore_388 replaced by KaratsubaCore_466

//KaratsubaCore_387 replaced by KaratsubaCore_465

//BADD_1589 replaced by BADD_1666

//BADD_1588 replaced by BADD_1668

//BADD_1587 replaced by BADD_1667

//BADD_1586 replaced by BADD_1666

//ADD_5487 replaced by ADD_8288

//ADD_5486 replaced by ADD_8288

//ADD_5485 replaced by ADD_8288

//ADD_5484 replaced by ADD_8288

//KaratsubaCore_392 replaced by KaratsubaCore_464

//KaratsubaCore_391 replaced by KaratsubaCore_463

//KaratsubaCore_390 replaced by KaratsubaCore_462

//BADD_1592 replaced by BADD_1672

//BADD_1591 replaced by BADD_1671

//BADD_1590 replaced by BADD_1670

//ADD_5491 replaced by ADD_11602

//ADD_5490 replaced by ADD_11602

//ADD_5489 replaced by ADD_11602

//ADD_5488 replaced by ADD_11602

//KaratsubaCore_395 replaced by KaratsubaCore_467

//KaratsubaCore_394 replaced by KaratsubaCore_466

//KaratsubaCore_393 replaced by KaratsubaCore_465

//ADD_5497 replaced by ADD_5761

//ADD_5496 replaced by ADD_5756

//ADD_5495 replaced by ADD_5756

//ADD_5494 replaced by ADD_5756

//ADD_5493 replaced by ADD_5756

//ADD_5492 replaced by ADD_5756

//ADD_5509 replaced by ADD_11602

//ADD_5508 replaced by ADD_11602

//ADD_5507 replaced by ADD_11602

//ADD_5506 replaced by ADD_11602

//ADD_5505 replaced by ADD_11602

//ADD_5504 replaced by ADD_11602

//ADD_5503 replaced by ADD_11602

//ADD_5502 replaced by ADD_11602

//ADD_5501 replaced by ADD_11602

//ADD_5500 replaced by ADD_11602

//ADD_5499 replaced by ADD_11602

//ADD_5498 replaced by ADD_11602

//ADD_5518 replaced by ADD_11601

//ADD_5517 replaced by ADD_11602

//ADD_5516 replaced by ADD_11602

//ADD_5515 replaced by ADD_11602

//ADD_5514 replaced by ADD_11602

//ADD_5513 replaced by ADD_11602

//ADD_5512 replaced by ADD_11602

//ADD_5511 replaced by ADD_11602

//ADD_5510 replaced by ADD_11602

//ADD_5526 replaced by ADD_11602

//ADD_5525 replaced by ADD_11602

//ADD_5524 replaced by ADD_11602

//ADD_5523 replaced by ADD_11602

//ADD_5522 replaced by ADD_11602

//ADD_5521 replaced by ADD_11602

//ADD_5520 replaced by ADD_11602

//ADD_5519 replaced by ADD_11602

//BADD_1595 replaced by BADD_1672

//BADD_1594 replaced by BADD_1671

//BADD_1593 replaced by BADD_1670

//ADD_5530 replaced by ADD_11602

//ADD_5529 replaced by ADD_11602

//ADD_5528 replaced by ADD_11602

//ADD_5527 replaced by ADD_11602

//KaratsubaCore_398 replaced by KaratsubaCore_467

//KaratsubaCore_397 replaced by KaratsubaCore_466

//KaratsubaCore_396 replaced by KaratsubaCore_465

//BADD_1599 replaced by BADD_1666

//BADD_1598 replaced by BADD_1668

//BADD_1597 replaced by BADD_1667

//BADD_1596 replaced by BADD_1666

//ADD_5534 replaced by ADD_8288

//ADD_5533 replaced by ADD_8288

//ADD_5532 replaced by ADD_8288

//ADD_5531 replaced by ADD_8288

//KaratsubaCore_401 replaced by KaratsubaCore_464

//KaratsubaCore_400 replaced by KaratsubaCore_463

//KaratsubaCore_399 replaced by KaratsubaCore_462

//BADD_1602 replaced by BADD_1672

//BADD_1601 replaced by BADD_1671

//BADD_1600 replaced by BADD_1670

//ADD_5538 replaced by ADD_11602

//ADD_5537 replaced by ADD_11602

//ADD_5536 replaced by ADD_11602

//ADD_5535 replaced by ADD_11602

//KaratsubaCore_404 replaced by KaratsubaCore_467

//KaratsubaCore_403 replaced by KaratsubaCore_466

//KaratsubaCore_402 replaced by KaratsubaCore_465

//ADD_5550 replaced by ADD_11602

//ADD_5549 replaced by ADD_11602

//ADD_5548 replaced by ADD_11602

//ADD_5547 replaced by ADD_11602

//ADD_5546 replaced by ADD_11602

//ADD_5545 replaced by ADD_11602

//ADD_5544 replaced by ADD_11602

//ADD_5543 replaced by ADD_11602

//ADD_5542 replaced by ADD_11602

//ADD_5541 replaced by ADD_11602

//ADD_5540 replaced by ADD_11602

//ADD_5539 replaced by ADD_11602

//ADD_5559 replaced by ADD_11601

//ADD_5558 replaced by ADD_11602

//ADD_5557 replaced by ADD_11602

//ADD_5556 replaced by ADD_11602

//ADD_5555 replaced by ADD_11602

//ADD_5554 replaced by ADD_11602

//ADD_5553 replaced by ADD_11602

//ADD_5552 replaced by ADD_11602

//ADD_5551 replaced by ADD_11602

//ADD_5567 replaced by ADD_11602

//ADD_5566 replaced by ADD_11602

//ADD_5565 replaced by ADD_11602

//ADD_5564 replaced by ADD_11602

//ADD_5563 replaced by ADD_11602

//ADD_5562 replaced by ADD_11602

//ADD_5561 replaced by ADD_11602

//ADD_5560 replaced by ADD_11602

//BADD_1605 replaced by BADD_1672

//BADD_1604 replaced by BADD_1671

//BADD_1603 replaced by BADD_1670

//ADD_5571 replaced by ADD_11602

//ADD_5570 replaced by ADD_11602

//ADD_5569 replaced by ADD_11602

//ADD_5568 replaced by ADD_11602

//KaratsubaCore_407 replaced by KaratsubaCore_467

//KaratsubaCore_406 replaced by KaratsubaCore_466

//KaratsubaCore_405 replaced by KaratsubaCore_465

//BADD_1609 replaced by BADD_1666

//BADD_1608 replaced by BADD_1668

//BADD_1607 replaced by BADD_1667

//BADD_1606 replaced by BADD_1666

//ADD_5575 replaced by ADD_8288

//ADD_5574 replaced by ADD_8288

//ADD_5573 replaced by ADD_8288

//ADD_5572 replaced by ADD_8288

//KaratsubaCore_410 replaced by KaratsubaCore_464

//KaratsubaCore_409 replaced by KaratsubaCore_463

//KaratsubaCore_408 replaced by KaratsubaCore_462

//BADD_1612 replaced by BADD_1672

//BADD_1611 replaced by BADD_1671

//BADD_1610 replaced by BADD_1670

//ADD_5579 replaced by ADD_11602

//ADD_5578 replaced by ADD_11602

//ADD_5577 replaced by ADD_11602

//ADD_5576 replaced by ADD_11602

//KaratsubaCore_413 replaced by KaratsubaCore_467

//KaratsubaCore_412 replaced by KaratsubaCore_466

//KaratsubaCore_411 replaced by KaratsubaCore_465

//ADD_5585 replaced by ADD_5761

//ADD_5584 replaced by ADD_5756

//ADD_5583 replaced by ADD_5756

//ADD_5582 replaced by ADD_5756

//ADD_5581 replaced by ADD_5756

//ADD_5580 replaced by ADD_5756

//ADD_5597 replaced by ADD_11602

//ADD_5596 replaced by ADD_11602

//ADD_5595 replaced by ADD_11602

//ADD_5594 replaced by ADD_11602

//ADD_5593 replaced by ADD_11602

//ADD_5592 replaced by ADD_11602

//ADD_5591 replaced by ADD_11602

//ADD_5590 replaced by ADD_11602

//ADD_5589 replaced by ADD_11602

//ADD_5588 replaced by ADD_11602

//ADD_5587 replaced by ADD_11602

//ADD_5586 replaced by ADD_11602

//ADD_5606 replaced by ADD_11601

//ADD_5605 replaced by ADD_11602

//ADD_5604 replaced by ADD_11602

//ADD_5603 replaced by ADD_11602

//ADD_5602 replaced by ADD_11602

//ADD_5601 replaced by ADD_11602

//ADD_5600 replaced by ADD_11602

//ADD_5599 replaced by ADD_11602

//ADD_5598 replaced by ADD_11602

//ADD_5614 replaced by ADD_11602

//ADD_5613 replaced by ADD_11602

//ADD_5612 replaced by ADD_11602

//ADD_5611 replaced by ADD_11602

//ADD_5610 replaced by ADD_11602

//ADD_5609 replaced by ADD_11602

//ADD_5608 replaced by ADD_11602

//ADD_5607 replaced by ADD_11602

//BADD_1615 replaced by BADD_1672

//BADD_1614 replaced by BADD_1671

//BADD_1613 replaced by BADD_1670

//ADD_5618 replaced by ADD_11602

//ADD_5617 replaced by ADD_11602

//ADD_5616 replaced by ADD_11602

//ADD_5615 replaced by ADD_11602

//KaratsubaCore_416 replaced by KaratsubaCore_467

//KaratsubaCore_415 replaced by KaratsubaCore_466

//KaratsubaCore_414 replaced by KaratsubaCore_465

//BADD_1619 replaced by BADD_1666

//BADD_1618 replaced by BADD_1668

//BADD_1617 replaced by BADD_1667

//BADD_1616 replaced by BADD_1666

//ADD_5622 replaced by ADD_8288

//ADD_5621 replaced by ADD_8288

//ADD_5620 replaced by ADD_8288

//ADD_5619 replaced by ADD_8288

//KaratsubaCore_419 replaced by KaratsubaCore_464

//KaratsubaCore_418 replaced by KaratsubaCore_463

//KaratsubaCore_417 replaced by KaratsubaCore_462

//BADD_1622 replaced by BADD_1672

//BADD_1621 replaced by BADD_1671

//BADD_1620 replaced by BADD_1670

//ADD_5626 replaced by ADD_11602

//ADD_5625 replaced by ADD_11602

//ADD_5624 replaced by ADD_11602

//ADD_5623 replaced by ADD_11602

//KaratsubaCore_422 replaced by KaratsubaCore_467

//KaratsubaCore_421 replaced by KaratsubaCore_466

//KaratsubaCore_420 replaced by KaratsubaCore_465

//ADD_5638 replaced by ADD_11602

//ADD_5637 replaced by ADD_11602

//ADD_5636 replaced by ADD_11602

//ADD_5635 replaced by ADD_11602

//ADD_5634 replaced by ADD_11602

//ADD_5633 replaced by ADD_11602

//ADD_5632 replaced by ADD_11602

//ADD_5631 replaced by ADD_11602

//ADD_5630 replaced by ADD_11602

//ADD_5629 replaced by ADD_11602

//ADD_5628 replaced by ADD_11602

//ADD_5627 replaced by ADD_11602

//ADD_5647 replaced by ADD_11601

//ADD_5646 replaced by ADD_11602

//ADD_5645 replaced by ADD_11602

//ADD_5644 replaced by ADD_11602

//ADD_5643 replaced by ADD_11602

//ADD_5642 replaced by ADD_11602

//ADD_5641 replaced by ADD_11602

//ADD_5640 replaced by ADD_11602

//ADD_5639 replaced by ADD_11602

//ADD_5655 replaced by ADD_11602

//ADD_5654 replaced by ADD_11602

//ADD_5653 replaced by ADD_11602

//ADD_5652 replaced by ADD_11602

//ADD_5651 replaced by ADD_11602

//ADD_5650 replaced by ADD_11602

//ADD_5649 replaced by ADD_11602

//ADD_5648 replaced by ADD_11602

//BADD_1625 replaced by BADD_1672

//BADD_1624 replaced by BADD_1671

//BADD_1623 replaced by BADD_1670

//ADD_5659 replaced by ADD_11602

//ADD_5658 replaced by ADD_11602

//ADD_5657 replaced by ADD_11602

//ADD_5656 replaced by ADD_11602

//KaratsubaCore_425 replaced by KaratsubaCore_467

//KaratsubaCore_424 replaced by KaratsubaCore_466

//KaratsubaCore_423 replaced by KaratsubaCore_465

//BADD_1629 replaced by BADD_1666

//BADD_1628 replaced by BADD_1668

//BADD_1627 replaced by BADD_1667

//BADD_1626 replaced by BADD_1666

//ADD_5663 replaced by ADD_8288

//ADD_5662 replaced by ADD_8288

//ADD_5661 replaced by ADD_8288

//ADD_5660 replaced by ADD_8288

//KaratsubaCore_428 replaced by KaratsubaCore_464

//KaratsubaCore_427 replaced by KaratsubaCore_463

//KaratsubaCore_426 replaced by KaratsubaCore_462

//BADD_1632 replaced by BADD_1672

//BADD_1631 replaced by BADD_1671

//BADD_1630 replaced by BADD_1670

//ADD_5667 replaced by ADD_11602

//ADD_5666 replaced by ADD_11602

//ADD_5665 replaced by ADD_11602

//ADD_5664 replaced by ADD_11602

//KaratsubaCore_431 replaced by KaratsubaCore_467

//KaratsubaCore_430 replaced by KaratsubaCore_466

//KaratsubaCore_429 replaced by KaratsubaCore_465

//ADD_5673 replaced by ADD_5761

//ADD_5672 replaced by ADD_5756

//ADD_5671 replaced by ADD_5756

//ADD_5670 replaced by ADD_5756

//ADD_5669 replaced by ADD_5756

//ADD_5668 replaced by ADD_5756

//ADD_5685 replaced by ADD_11602

//ADD_5684 replaced by ADD_11602

//ADD_5683 replaced by ADD_11602

//ADD_5682 replaced by ADD_11602

//ADD_5681 replaced by ADD_11602

//ADD_5680 replaced by ADD_11602

//ADD_5679 replaced by ADD_11602

//ADD_5678 replaced by ADD_11602

//ADD_5677 replaced by ADD_11602

//ADD_5676 replaced by ADD_11602

//ADD_5675 replaced by ADD_11602

//ADD_5674 replaced by ADD_11602

//ADD_5694 replaced by ADD_11601

//ADD_5693 replaced by ADD_11602

//ADD_5692 replaced by ADD_11602

//ADD_5691 replaced by ADD_11602

//ADD_5690 replaced by ADD_11602

//ADD_5689 replaced by ADD_11602

//ADD_5688 replaced by ADD_11602

//ADD_5687 replaced by ADD_11602

//ADD_5686 replaced by ADD_11602

//ADD_5702 replaced by ADD_11602

//ADD_5701 replaced by ADD_11602

//ADD_5700 replaced by ADD_11602

//ADD_5699 replaced by ADD_11602

//ADD_5698 replaced by ADD_11602

//ADD_5697 replaced by ADD_11602

//ADD_5696 replaced by ADD_11602

//ADD_5695 replaced by ADD_11602

//BADD_1635 replaced by BADD_1672

//BADD_1634 replaced by BADD_1671

//BADD_1633 replaced by BADD_1670

//ADD_5706 replaced by ADD_11602

//ADD_5705 replaced by ADD_11602

//ADD_5704 replaced by ADD_11602

//ADD_5703 replaced by ADD_11602

//KaratsubaCore_434 replaced by KaratsubaCore_467

//KaratsubaCore_433 replaced by KaratsubaCore_466

//KaratsubaCore_432 replaced by KaratsubaCore_465

//BADD_1639 replaced by BADD_1666

//BADD_1638 replaced by BADD_1668

//BADD_1637 replaced by BADD_1667

//BADD_1636 replaced by BADD_1666

//ADD_5710 replaced by ADD_8288

//ADD_5709 replaced by ADD_8288

//ADD_5708 replaced by ADD_8288

//ADD_5707 replaced by ADD_8288

//KaratsubaCore_437 replaced by KaratsubaCore_464

//KaratsubaCore_436 replaced by KaratsubaCore_463

//KaratsubaCore_435 replaced by KaratsubaCore_462

//BADD_1642 replaced by BADD_1672

//BADD_1641 replaced by BADD_1671

//BADD_1640 replaced by BADD_1670

//ADD_5714 replaced by ADD_11602

//ADD_5713 replaced by ADD_11602

//ADD_5712 replaced by ADD_11602

//ADD_5711 replaced by ADD_11602

//KaratsubaCore_440 replaced by KaratsubaCore_467

//KaratsubaCore_439 replaced by KaratsubaCore_466

//KaratsubaCore_438 replaced by KaratsubaCore_465

//ADD_5726 replaced by ADD_11602

//ADD_5725 replaced by ADD_11602

//ADD_5724 replaced by ADD_11602

//ADD_5723 replaced by ADD_11602

//ADD_5722 replaced by ADD_11602

//ADD_5721 replaced by ADD_11602

//ADD_5720 replaced by ADD_11602

//ADD_5719 replaced by ADD_11602

//ADD_5718 replaced by ADD_11602

//ADD_5717 replaced by ADD_11602

//ADD_5716 replaced by ADD_11602

//ADD_5715 replaced by ADD_11602

//ADD_5735 replaced by ADD_11601

//ADD_5734 replaced by ADD_11602

//ADD_5733 replaced by ADD_11602

//ADD_5732 replaced by ADD_11602

//ADD_5731 replaced by ADD_11602

//ADD_5730 replaced by ADD_11602

//ADD_5729 replaced by ADD_11602

//ADD_5728 replaced by ADD_11602

//ADD_5727 replaced by ADD_11602

//ADD_5743 replaced by ADD_11602

//ADD_5742 replaced by ADD_11602

//ADD_5741 replaced by ADD_11602

//ADD_5740 replaced by ADD_11602

//ADD_5739 replaced by ADD_11602

//ADD_5738 replaced by ADD_11602

//ADD_5737 replaced by ADD_11602

//ADD_5736 replaced by ADD_11602

//BADD_1645 replaced by BADD_1672

//BADD_1644 replaced by BADD_1671

//BADD_1643 replaced by BADD_1670

//ADD_5747 replaced by ADD_11602

//ADD_5746 replaced by ADD_11602

//ADD_5745 replaced by ADD_11602

//ADD_5744 replaced by ADD_11602

//KaratsubaCore_443 replaced by KaratsubaCore_467

//KaratsubaCore_442 replaced by KaratsubaCore_466

//KaratsubaCore_441 replaced by KaratsubaCore_465

//BADD_1649 replaced by BADD_1666

//BADD_1648 replaced by BADD_1668

//BADD_1647 replaced by BADD_1667

//BADD_1646 replaced by BADD_1666

//ADD_5751 replaced by ADD_8288

//ADD_5750 replaced by ADD_8288

//ADD_5749 replaced by ADD_8288

//ADD_5748 replaced by ADD_8288

//KaratsubaCore_446 replaced by KaratsubaCore_464

//KaratsubaCore_445 replaced by KaratsubaCore_463

//KaratsubaCore_444 replaced by KaratsubaCore_462

//BADD_1652 replaced by BADD_1672

//BADD_1651 replaced by BADD_1671

//BADD_1650 replaced by BADD_1670

//ADD_5755 replaced by ADD_11602

//ADD_5754 replaced by ADD_11602

//ADD_5753 replaced by ADD_11602

//ADD_5752 replaced by ADD_11602

//KaratsubaCore_449 replaced by KaratsubaCore_467

//KaratsubaCore_448 replaced by KaratsubaCore_466

//KaratsubaCore_447 replaced by KaratsubaCore_465

module ADD_5761 (
  input      [57:0]   io_A_0,
  input      [57:0]   io_A_1,
  input               io_CIN,
  output     [58:0]   io_S
);

  wire       [58:0]   _zz_io_S;
  wire       [58:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {58'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_5760 replaced by ADD_5756

//ADD_5759 replaced by ADD_5756

//ADD_5758 replaced by ADD_5756

//ADD_5757 replaced by ADD_5756

module ADD_5756 (
  input      [63:0]   io_A_0,
  input      [63:0]   io_A_1,
  input               io_CIN,
  output     [64:0]   io_S
);

  wire       [64:0]   _zz_io_S;
  wire       [64:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {64'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_5773 replaced by ADD_11602

//ADD_5772 replaced by ADD_11602

//ADD_5771 replaced by ADD_11602

//ADD_5770 replaced by ADD_11602

//ADD_5769 replaced by ADD_11602

//ADD_5768 replaced by ADD_11602

//ADD_5767 replaced by ADD_11602

//ADD_5766 replaced by ADD_11602

//ADD_5765 replaced by ADD_11602

//ADD_5764 replaced by ADD_11602

//ADD_5763 replaced by ADD_11602

//ADD_5762 replaced by ADD_11602

//ADD_5782 replaced by ADD_11601

//ADD_5781 replaced by ADD_11602

//ADD_5780 replaced by ADD_11602

//ADD_5779 replaced by ADD_11602

//ADD_5778 replaced by ADD_11602

//ADD_5777 replaced by ADD_11602

//ADD_5776 replaced by ADD_11602

//ADD_5775 replaced by ADD_11602

//ADD_5774 replaced by ADD_11602

//ADD_5790 replaced by ADD_11602

//ADD_5789 replaced by ADD_11602

//ADD_5788 replaced by ADD_11602

//ADD_5787 replaced by ADD_11602

//ADD_5786 replaced by ADD_11602

//ADD_5785 replaced by ADD_11602

//ADD_5784 replaced by ADD_11602

//ADD_5783 replaced by ADD_11602

//BADD_1655 replaced by BADD_1672

//BADD_1654 replaced by BADD_1671

//BADD_1653 replaced by BADD_1670

//ADD_5794 replaced by ADD_11602

//ADD_5793 replaced by ADD_11602

//ADD_5792 replaced by ADD_11602

//ADD_5791 replaced by ADD_11602

//KaratsubaCore_452 replaced by KaratsubaCore_467

//KaratsubaCore_451 replaced by KaratsubaCore_466

//KaratsubaCore_450 replaced by KaratsubaCore_465

//BADD_1659 replaced by BADD_1666

//BADD_1658 replaced by BADD_1668

//BADD_1657 replaced by BADD_1667

//BADD_1656 replaced by BADD_1666

//ADD_5798 replaced by ADD_8288

//ADD_5797 replaced by ADD_8288

//ADD_5796 replaced by ADD_8288

//ADD_5795 replaced by ADD_8288

//KaratsubaCore_455 replaced by KaratsubaCore_464

//KaratsubaCore_454 replaced by KaratsubaCore_463

//KaratsubaCore_453 replaced by KaratsubaCore_462

//BADD_1662 replaced by BADD_1672

//BADD_1661 replaced by BADD_1671

//BADD_1660 replaced by BADD_1670

//ADD_5802 replaced by ADD_11602

//ADD_5801 replaced by ADD_11602

//ADD_5800 replaced by ADD_11602

//ADD_5799 replaced by ADD_11602

//KaratsubaCore_458 replaced by KaratsubaCore_467

//KaratsubaCore_457 replaced by KaratsubaCore_466

//KaratsubaCore_456 replaced by KaratsubaCore_465

//ADD_5814 replaced by ADD_11602

//ADD_5813 replaced by ADD_11602

//ADD_5812 replaced by ADD_11602

//ADD_5811 replaced by ADD_11602

//ADD_5810 replaced by ADD_11602

//ADD_5809 replaced by ADD_11602

//ADD_5808 replaced by ADD_11602

//ADD_5807 replaced by ADD_11602

//ADD_5806 replaced by ADD_11602

//ADD_5805 replaced by ADD_11602

//ADD_5804 replaced by ADD_11602

//ADD_5803 replaced by ADD_11602

//ADD_5823 replaced by ADD_11601

//ADD_5822 replaced by ADD_11602

//ADD_5821 replaced by ADD_11602

//ADD_5820 replaced by ADD_11602

//ADD_5819 replaced by ADD_11602

//ADD_5818 replaced by ADD_11602

//ADD_5817 replaced by ADD_11602

//ADD_5816 replaced by ADD_11602

//ADD_5815 replaced by ADD_11602

//ADD_5831 replaced by ADD_11602

//ADD_5830 replaced by ADD_11602

//ADD_5829 replaced by ADD_11602

//ADD_5828 replaced by ADD_11602

//ADD_5827 replaced by ADD_11602

//ADD_5826 replaced by ADD_11602

//ADD_5825 replaced by ADD_11602

//ADD_5824 replaced by ADD_11602

//BADD_1665 replaced by BADD_1672

//BADD_1664 replaced by BADD_1671

//BADD_1663 replaced by BADD_1670

//ADD_5835 replaced by ADD_11602

//ADD_5834 replaced by ADD_11602

//ADD_5833 replaced by ADD_11602

//ADD_5832 replaced by ADD_11602

//KaratsubaCore_461 replaced by KaratsubaCore_467

//KaratsubaCore_460 replaced by KaratsubaCore_466

//KaratsubaCore_459 replaced by KaratsubaCore_465

//BADD_1669 replaced by BADD_1666

module BADD_1668 (
  input      [194:0]  io_a,
  input      [194:0]  io_b,
  input               io_c,
  output     [195:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [2:0]    adder_adds_4_io_A_0;
  wire       [2:0]    adder_adds_4_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  wire       [3:0]    adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [2:0]    _zz_io_s_5;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  ADD_11592 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[2:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[2:0]), //i
    .io_CIN (_zz_io_CIN_3            ), //i
    .io_S   (adder_adds_4_io_S[3:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_4_io_A_0 = io_a[194 : 192];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[143 : 96];
  assign adder_adds_3_io_A_1 = io_b[191 : 144];
  assign adder_adds_4_io_A_1 = io_b[194 : 192];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_CIN_3 <= adder_adds_3_io_S[48];
    _zz_io_s <= adder_adds_4_io_S[3];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[2 : 0];
  end


endmodule

module BADD_1667 (
  input      [194:0]  io_a,
  input      [194:0]  io_b,
  input               io_c,
  output     [195:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [2:0]    adder_adds_4_io_A_0;
  wire       [2:0]    adder_adds_4_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  wire       [3:0]    adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [2:0]    _zz_io_s_5;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  ADD_11592 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[2:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[2:0]), //i
    .io_CIN (_zz_io_CIN_3            ), //i
    .io_S   (adder_adds_4_io_S[3:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_4_io_A_0 = io_a[194 : 192];
  assign adder_adds_0_io_A_1 = (~ io_b[47 : 0]);
  assign adder_adds_1_io_A_1 = (~ io_b[95 : 48]);
  assign adder_adds_2_io_A_1 = (~ io_b[143 : 96]);
  assign adder_adds_3_io_A_1 = (~ io_b[191 : 144]);
  assign adder_adds_4_io_A_1 = (~ io_b[194 : 192]);
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_CIN_3 <= adder_adds_3_io_S[48];
    _zz_io_s <= (! adder_adds_4_io_S[3]);
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[2 : 0];
  end


endmodule

module BADD_1666 (
  input      [193:0]  io_a,
  input      [193:0]  io_b,
  input               io_c,
  output     [194:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [1:0]    adder_adds_4_io_A_0;
  wire       [1:0]    adder_adds_4_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  wire       [2:0]    adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [1:0]    _zz_io_s_5;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  ADD_11595 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[1:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[1:0]), //i
    .io_CIN (_zz_io_CIN_3            ), //i
    .io_S   (adder_adds_4_io_S[2:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_4_io_A_0 = io_a[193 : 192];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[143 : 96];
  assign adder_adds_3_io_A_1 = io_b[191 : 144];
  assign adder_adds_4_io_A_1 = io_b[193 : 192];
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_CIN_3 <= adder_adds_3_io_S[48];
    _zz_io_s <= adder_adds_4_io_S[2];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[1 : 0];
  end


endmodule

//ADD_5839 replaced by ADD_8288

//ADD_5838 replaced by ADD_8288

//ADD_5837 replaced by ADD_8288

//ADD_5836 replaced by ADD_8288

module KaratsubaCore_464 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_a_1,
  input      [48:0]   io_b_0,
  input      [48:0]   io_b_1,
  output reg [193:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [98:0]   karatsuba_add2_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_b;
  wire       [97:0]   karatsuba_hasExtend_add4_io_a;
  wire       [97:0]   karatsuba_lsbMul_io_p;
  wire       [99:0]   karatsuba_midMul_io_p;
  wire       [97:0]   karatsuba_msbMul_io_p;
  wire       [49:0]   karatsuba_midAdd_0_0_io_S;
  wire       [49:0]   karatsuba_midAdd_1_0_io_S;
  wire       [98:0]   karatsuba_add1_io_s;
  wire       [99:0]   karatsuba_add2_io_s;
  wire       [99:0]   karatsuba_hasExtend_add3_io_s;
  wire       [98:0]   karatsuba_hasExtend_add4_io_s;
  wire       [51:0]   _zz_io_a;
  reg        [49:0]   _zz_io_a_0;
  reg        [49:0]   _zz_io_b_0;
  reg        [49:0]   _zz_io_b;
  reg        [97:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [97:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [97:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [97:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;

  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 48);
  KaratsubaCore_1438 karatsuba_lsbMul (
    .io_a_0 (io_a_0[48:0]               ), //i
    .io_b_0 (io_b_0[48:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1435 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[49:0]           ), //i
    .io_b_0 (_zz_io_b_0[49:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1438 karatsuba_msbMul (
    .io_a_0 (io_a_1[48:0]               ), //i
    .io_b_0 (io_b_1[48:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  ADD_8288 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[48:0]                   ), //i
    .io_A_1 (io_a_1[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[49:0])  //o
  );
  ADD_8288 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[48:0]                   ), //i
    .io_A_1 (io_b_1[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[49:0])  //o
  );
  BADD_2818 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[97:0]), //i
    .io_b   (karatsuba_msbMul_io_p[97:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[98:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_2819 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[98:0]), //i
    .io_b   (karatsuba_add1_io_s[98:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[99:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_2820 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[98:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[98:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[99:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  BADD_2818 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[97:0]                 ), //i
    .io_b   (karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4[97:0]), //i
    .io_c   (1'b0                                                ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[98:0]                 ), //o
    .clk    (clk                                                 ), //i
    .resetn (resetn                                              )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[98:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[98:0];
  assign karatsuba_hasExtend_add3_io_b = {49'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {46'd0, _zz_io_a};
  always @(*) begin
    io_p[47 : 0] = _zz_io_p_2;
    io_p[95 : 48] = _zz_io_p_3;
    io_p[193 : 96] = karatsuba_hasExtend_add4_io_s[97:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= karatsuba_hasExtend_add3_io_s[47:0];
  end


endmodule

module KaratsubaCore_463 (
  input      [49:0]   io_a_0,
  input      [49:0]   io_a_1,
  input      [49:0]   io_b_0,
  input      [49:0]   io_b_1,
  output reg [195:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [100:0]  karatsuba_add2_io_a;
  wire       [100:0]  karatsuba_hasExtend_add3_io_a;
  wire       [100:0]  karatsuba_hasExtend_add3_io_b;
  wire       [99:0]   karatsuba_hasExtend_add4_io_a;
  wire       [99:0]   karatsuba_lsbMul_io_p;
  wire       [101:0]  karatsuba_midMul_io_p;
  wire       [99:0]   karatsuba_msbMul_io_p;
  wire       [50:0]   karatsuba_midAdd_0_0_io_S;
  wire       [50:0]   karatsuba_midAdd_1_0_io_S;
  wire       [100:0]  karatsuba_add1_io_s;
  wire       [101:0]  karatsuba_add2_io_s;
  wire       [101:0]  karatsuba_hasExtend_add3_io_s;
  wire       [100:0]  karatsuba_hasExtend_add4_io_s;
  wire       [53:0]   _zz_io_a;
  reg        [50:0]   _zz_io_a_0;
  reg        [50:0]   _zz_io_b_0;
  reg        [51:0]   _zz_io_b;
  reg        [99:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
  reg        [99:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
  reg        [99:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
  reg        [99:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_4;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;

  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 48);
  KaratsubaCore_1435 karatsuba_lsbMul (
    .io_a_0 (io_a_0[49:0]               ), //i
    .io_b_0 (io_b_0[49:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1426 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[50:0]            ), //i
    .io_b_0 (_zz_io_b_0[50:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[101:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_1435 karatsuba_msbMul (
    .io_a_0 (io_a_1[49:0]               ), //i
    .io_b_0 (io_b_1[49:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  ADD_8267 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[49:0]                   ), //i
    .io_A_1 (io_a_1[49:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[50:0])  //o
  );
  ADD_8267 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[49:0]                   ), //i
    .io_A_1 (io_b_1[49:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[50:0])  //o
  );
  BADD_2807 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[99:0]), //i
    .io_b   (karatsuba_msbMul_io_p[99:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[100:0] ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_2808 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[100:0]), //i
    .io_b   (karatsuba_add1_io_s[100:0]), //i
    .io_c   (1'b1                      ), //i
    .io_s   (karatsuba_add2_io_s[101:0]), //o
    .clk    (clk                       ), //i
    .resetn (resetn                    )  //i
  );
  BADD_2809 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[100:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[100:0]), //i
    .io_c   (1'b0                                ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[101:0]), //o
    .clk    (clk                                 ), //i
    .resetn (resetn                              )  //i
  );
  BADD_2807 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[99:0]                 ), //i
    .io_b   (karatsuba_midMul_karatsuba_msbMul_io_p_delay_4[99:0]), //i
    .io_c   (1'b0                                                ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[100:0]                ), //o
    .clk    (clk                                                 ), //i
    .resetn (resetn                                              )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[100:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[100:0];
  assign karatsuba_hasExtend_add3_io_b = {49'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {46'd0, _zz_io_a};
  always @(*) begin
    io_p[47 : 0] = _zz_io_p_2;
    io_p[95 : 48] = _zz_io_p_3;
    io_p[195 : 96] = karatsuba_hasExtend_add4_io_s[99:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= karatsuba_hasExtend_add3_io_s[47:0];
  end


endmodule

module KaratsubaCore_462 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_a_1,
  input      [48:0]   io_b_0,
  input      [48:0]   io_b_1,
  output reg [193:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [98:0]   karatsuba_add2_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_b;
  wire       [97:0]   karatsuba_hasExtend_add4_io_a;
  wire       [97:0]   karatsuba_lsbMul_io_p;
  wire       [99:0]   karatsuba_midMul_io_p;
  wire       [97:0]   karatsuba_msbMul_io_p;
  wire       [49:0]   karatsuba_midAdd_0_0_io_S;
  wire       [49:0]   karatsuba_midAdd_1_0_io_S;
  wire       [98:0]   karatsuba_add1_io_s;
  wire       [99:0]   karatsuba_add2_io_s;
  wire       [99:0]   karatsuba_hasExtend_add3_io_s;
  wire       [98:0]   karatsuba_hasExtend_add4_io_s;
  wire       [51:0]   _zz_io_a;
  reg        [49:0]   _zz_io_a_0;
  reg        [49:0]   _zz_io_b_0;
  reg        [49:0]   _zz_io_b;
  reg        [97:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [97:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [97:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [97:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;

  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 48);
  KaratsubaCore_1438 karatsuba_lsbMul (
    .io_a_0 (io_a_0[48:0]               ), //i
    .io_b_0 (io_b_0[48:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1435 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[49:0]           ), //i
    .io_b_0 (_zz_io_b_0[49:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1438 karatsuba_msbMul (
    .io_a_0 (io_a_1[48:0]               ), //i
    .io_b_0 (io_b_1[48:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  ADD_8288 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[48:0]                   ), //i
    .io_A_1 (io_a_1[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[49:0])  //o
  );
  ADD_8288 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[48:0]                   ), //i
    .io_A_1 (io_b_1[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[49:0])  //o
  );
  BADD_2818 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[97:0]), //i
    .io_b   (karatsuba_msbMul_io_p[97:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[98:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_2819 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[98:0]), //i
    .io_b   (karatsuba_add1_io_s[98:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[99:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_2820 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[98:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[98:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[99:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  BADD_2818 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[97:0]                 ), //i
    .io_b   (karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4[97:0]), //i
    .io_c   (1'b0                                                ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[98:0]                 ), //o
    .clk    (clk                                                 ), //i
    .resetn (resetn                                              )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[98:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[98:0];
  assign karatsuba_hasExtend_add3_io_b = {49'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {46'd0, _zz_io_a};
  always @(*) begin
    io_p[47 : 0] = _zz_io_p_2;
    io_p[95 : 48] = _zz_io_p_3;
    io_p[193 : 96] = karatsuba_hasExtend_add4_io_s[97:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= karatsuba_hasExtend_add3_io_s[47:0];
  end


endmodule

module BADD_1672 (
  input      [287:0]  io_a,
  input      [287:0]  io_b,
  input               io_c,
  output     [288:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [47:0]   adder_adds_4_io_A_0;
  wire       [47:0]   adder_adds_4_io_A_1;
  wire       [47:0]   adder_adds_5_io_A_0;
  wire       [47:0]   adder_adds_5_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  wire       [48:0]   adder_adds_4_io_S;
  wire       [48:0]   adder_adds_5_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_CIN_4;
  reg                 _zz_io_s;
  reg                 _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [47:0]   _zz_io_s_5;
  reg        [47:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_4_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_3             ), //i
    .io_S   (adder_adds_4_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_5 (
    .io_A_0 (adder_adds_5_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_5_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_4             ), //i
    .io_S   (adder_adds_5_io_S[48:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_4_io_A_0 = io_a[239 : 192];
  assign adder_adds_5_io_A_0 = io_a[287 : 240];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[143 : 96];
  assign adder_adds_3_io_A_1 = io_b[191 : 144];
  assign adder_adds_4_io_A_1 = io_b[239 : 192];
  assign adder_adds_5_io_A_1 = io_b[287 : 240];
  assign io_s = {_zz_io_s_1,{_zz_io_s_7,{_zz_io_s_6,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,_zz_io_s_2}}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_CIN_3 <= adder_adds_3_io_S[48];
    _zz_io_CIN_4 <= adder_adds_4_io_S[48];
    _zz_io_s <= adder_adds_5_io_S[48];
    _zz_io_s_1 <= _zz_io_s;
    _zz_io_s_2 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_3_io_S[47 : 0];
    _zz_io_s_6 <= adder_adds_4_io_S[47 : 0];
    _zz_io_s_7 <= adder_adds_5_io_S[47 : 0];
  end


endmodule

module BADD_1671 (
  input      [192:0]  io_a,
  input      [192:0]  io_b,
  input               io_c,
  output     [193:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [0:0]    adder_adds_4_io_A_0;
  wire       [0:0]    adder_adds_4_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  wire       [1:0]    adder_adds_4_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_CIN_3;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [0:0]    _zz_io_s_5;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  ADD_11601 adder_adds_4 (
    .io_A_0 (adder_adds_4_io_A_0   ), //i
    .io_A_1 (adder_adds_4_io_A_1   ), //i
    .io_CIN (_zz_io_CIN_3          ), //i
    .io_S   (adder_adds_4_io_S[1:0])  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_4_io_A_0 = io_a[192 : 192];
  assign adder_adds_0_io_A_1 = (~ io_b[47 : 0]);
  assign adder_adds_1_io_A_1 = (~ io_b[95 : 48]);
  assign adder_adds_2_io_A_1 = (~ io_b[143 : 96]);
  assign adder_adds_3_io_A_1 = (~ io_b[191 : 144]);
  assign adder_adds_4_io_A_1 = (~ io_b[192 : 192]);
  assign io_s = {_zz_io_s,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_CIN_3 <= adder_adds_3_io_S[48];
    _zz_io_s <= (! adder_adds_4_io_S[1]);
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_3_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_4_io_S[0 : 0];
  end


endmodule

module BADD_1670 (
  input      [191:0]  io_a,
  input      [191:0]  io_b,
  input               io_c,
  output     [192:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [47:0]   adder_adds_3_io_A_0;
  wire       [47:0]   adder_adds_3_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  wire       [48:0]   adder_adds_3_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_CIN_2;
  reg                 _zz_io_s;
  reg                 _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg        [47:0]   _zz_io_s_5;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_3 (
    .io_A_0 (adder_adds_3_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_3_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_2             ), //i
    .io_S   (adder_adds_3_io_S[48:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_3_io_A_0 = io_a[191 : 144];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[143 : 96];
  assign adder_adds_3_io_A_1 = io_b[191 : 144];
  assign io_s = {_zz_io_s_1,{_zz_io_s_5,{_zz_io_s_4,{_zz_io_s_3,_zz_io_s_2}}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_CIN_2 <= adder_adds_2_io_S[48];
    _zz_io_s <= adder_adds_3_io_S[48];
    _zz_io_s_1 <= _zz_io_s;
    _zz_io_s_2 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_2_io_S[47 : 0];
    _zz_io_s_5 <= adder_adds_3_io_S[47 : 0];
  end


endmodule

//ADD_5843 replaced by ADD_11602

//ADD_5842 replaced by ADD_11602

//ADD_5841 replaced by ADD_11602

//ADD_5840 replaced by ADD_11602

module KaratsubaCore_467 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  output reg [191:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [96:0]   karatsuba_add2_io_a;
  wire       [143:0]  karatsuba_noExtend_add3_io_a;
  reg        [143:0]  karatsuba_noExtend_add3_io_b;
  wire       [95:0]   karatsuba_lsbMul_io_p;
  wire       [97:0]   karatsuba_midMul_io_p;
  wire       [95:0]   karatsuba_msbMul_io_p;
  wire       [48:0]   karatsuba_midAdd_0_0_io_S;
  wire       [48:0]   karatsuba_midAdd_1_0_io_S;
  wire       [96:0]   karatsuba_add1_io_s;
  wire       [97:0]   karatsuba_add2_io_s;
  wire       [144:0]  karatsuba_noExtend_add3_io_s;
  wire       [96:0]   _zz_io_a;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_b_0;
  reg        [47:0]   _zz_io_b;
  reg        [95:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [95:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [95:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;

  assign _zz_io_a = karatsuba_add2_io_s[96:0];
  KaratsubaCore_1437 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]               ), //i
    .io_b_0 (io_b_0[47:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[95:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1438 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]           ), //i
    .io_b_0 (_zz_io_b_0[48:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1437 karatsuba_msbMul (
    .io_a_0 (io_a_1[47:0]               ), //i
    .io_b_0 (io_b_1[47:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[95:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  ADD_11602 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[47:0]                   ), //i
    .io_A_1 (io_a_1[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[47:0]                   ), //i
    .io_A_1 (io_b_1[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[48:0])  //o
  );
  BADD_2822 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[95:0]), //i
    .io_b   (karatsuba_msbMul_io_p[95:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[96:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_2823 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[96:0]), //i
    .io_b   (karatsuba_add1_io_s[96:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[97:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_2824 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[143:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[143:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[144:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[96:0];
  assign karatsuba_noExtend_add3_io_a = {47'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[47 : 0] = _zz_io_b;
    karatsuba_noExtend_add3_io_b[143 : 48] = karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
  end

  always @(*) begin
    io_p[47 : 0] = _zz_io_p_1;
    io_p[191 : 48] = karatsuba_noExtend_add3_io_s[143:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
  end


endmodule

module KaratsubaCore_466 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_a_1,
  input      [48:0]   io_b_0,
  input      [48:0]   io_b_1,
  output reg [193:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [98:0]   karatsuba_add2_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_b;
  wire       [97:0]   karatsuba_hasExtend_add4_io_a;
  wire       [97:0]   karatsuba_lsbMul_io_p;
  wire       [99:0]   karatsuba_midMul_io_p;
  wire       [97:0]   karatsuba_msbMul_io_p;
  wire       [49:0]   karatsuba_midAdd_0_0_io_S;
  wire       [49:0]   karatsuba_midAdd_1_0_io_S;
  wire       [98:0]   karatsuba_add1_io_s;
  wire       [99:0]   karatsuba_add2_io_s;
  wire       [99:0]   karatsuba_hasExtend_add3_io_s;
  wire       [98:0]   karatsuba_hasExtend_add4_io_s;
  wire       [51:0]   _zz_io_a;
  reg        [49:0]   _zz_io_a_0;
  reg        [49:0]   _zz_io_b_0;
  reg        [49:0]   _zz_io_b;
  reg        [97:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
  reg        [97:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
  reg        [97:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
  reg        [97:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_4;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;

  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 48);
  KaratsubaCore_1438 karatsuba_lsbMul (
    .io_a_0 (io_a_0[48:0]               ), //i
    .io_b_0 (io_b_0[48:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1435 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[49:0]           ), //i
    .io_b_0 (_zz_io_b_0[49:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1438 karatsuba_msbMul (
    .io_a_0 (io_a_1[48:0]               ), //i
    .io_b_0 (io_b_1[48:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  ADD_8288 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[48:0]                   ), //i
    .io_A_1 (io_a_1[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[49:0])  //o
  );
  ADD_8288 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[48:0]                   ), //i
    .io_A_1 (io_b_1[48:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[49:0])  //o
  );
  BADD_2818 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[97:0]), //i
    .io_b   (karatsuba_msbMul_io_p[97:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[98:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_2819 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[98:0]), //i
    .io_b   (karatsuba_add1_io_s[98:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[99:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_2820 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[98:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[98:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[99:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  BADD_2818 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[97:0]                 ), //i
    .io_b   (karatsuba_midMul_karatsuba_msbMul_io_p_delay_4[97:0]), //i
    .io_c   (1'b0                                                ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[98:0]                 ), //o
    .clk    (clk                                                 ), //i
    .resetn (resetn                                              )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[98:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[98:0];
  assign karatsuba_hasExtend_add3_io_b = {49'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {46'd0, _zz_io_a};
  always @(*) begin
    io_p[47 : 0] = _zz_io_p_2;
    io_p[95 : 48] = _zz_io_p_3;
    io_p[193 : 96] = karatsuba_hasExtend_add4_io_s[97:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= karatsuba_hasExtend_add3_io_s[47:0];
  end


endmodule

module KaratsubaCore_465 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  output reg [191:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [96:0]   karatsuba_add2_io_a;
  wire       [143:0]  karatsuba_noExtend_add3_io_a;
  reg        [143:0]  karatsuba_noExtend_add3_io_b;
  wire       [95:0]   karatsuba_lsbMul_io_p;
  wire       [97:0]   karatsuba_midMul_io_p;
  wire       [95:0]   karatsuba_msbMul_io_p;
  wire       [48:0]   karatsuba_midAdd_0_0_io_S;
  wire       [48:0]   karatsuba_midAdd_1_0_io_S;
  wire       [96:0]   karatsuba_add1_io_s;
  wire       [97:0]   karatsuba_add2_io_s;
  wire       [144:0]  karatsuba_noExtend_add3_io_s;
  wire       [96:0]   _zz_io_a;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_b_0;
  reg        [47:0]   _zz_io_b;
  reg        [95:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [95:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [95:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;

  assign _zz_io_a = karatsuba_add2_io_s[96:0];
  KaratsubaCore_1437 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]               ), //i
    .io_b_0 (io_b_0[47:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[95:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1438 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]           ), //i
    .io_b_0 (_zz_io_b_0[48:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_1437 karatsuba_msbMul (
    .io_a_0 (io_a_1[47:0]               ), //i
    .io_b_0 (io_b_1[47:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[95:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  ADD_11602 karatsuba_midAdd_0_0 (
    .io_A_0 (io_a_0[47:0]                   ), //i
    .io_A_1 (io_a_1[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_0_0_io_S[48:0])  //o
  );
  ADD_11602 karatsuba_midAdd_1_0 (
    .io_A_0 (io_b_0[47:0]                   ), //i
    .io_A_1 (io_b_1[47:0]                   ), //i
    .io_CIN (1'b0                           ), //i
    .io_S   (karatsuba_midAdd_1_0_io_S[48:0])  //o
  );
  BADD_2822 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[95:0]), //i
    .io_b   (karatsuba_msbMul_io_p[95:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[96:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_2823 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[96:0]), //i
    .io_b   (karatsuba_add1_io_s[96:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[97:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_2824 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[143:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[143:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[144:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[96:0];
  assign karatsuba_noExtend_add3_io_a = {47'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[47 : 0] = _zz_io_b;
    karatsuba_noExtend_add3_io_b[143 : 48] = karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
  end

  always @(*) begin
    io_p[47 : 0] = _zz_io_p_1;
    io_p[191 : 48] = karatsuba_noExtend_add3_io_s[143:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= karatsuba_midAdd_0_0_io_S;
    _zz_io_b_0 <= karatsuba_midAdd_1_0_io_S;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
  end


endmodule

//ADD_5849 replaced by ADD_11602

//ADD_5848 replaced by ADD_11602

//ADD_5847 replaced by ADD_11602

//ADD_5846 replaced by ADD_11602

//ADD_5845 replaced by ADD_11602

//ADD_5844 replaced by ADD_11602

//ADD_5854 replaced by ADD_11601

//ADD_5853 replaced by ADD_11602

//ADD_5852 replaced by ADD_11602

//ADD_5851 replaced by ADD_11602

//ADD_5850 replaced by ADD_11602

//ADD_5858 replaced by ADD_11602

//ADD_5857 replaced by ADD_11602

//ADD_5856 replaced by ADD_11602

//ADD_5855 replaced by ADD_11602

//BADD_1675 replaced by BADD_2824

//BADD_1674 replaced by BADD_2823

//BADD_1673 replaced by BADD_2822

//ADD_5860 replaced by ADD_11602

//ADD_5859 replaced by ADD_11602

//KaratsubaCore_470 replaced by KaratsubaCore_1437

//KaratsubaCore_469 replaced by KaratsubaCore_1438

//KaratsubaCore_468 replaced by KaratsubaCore_1437

//BADD_1679 replaced by BADD_2818

//BADD_1678 replaced by BADD_2820

//BADD_1677 replaced by BADD_2819

//BADD_1676 replaced by BADD_2818

//ADD_5862 replaced by ADD_8288

//ADD_5861 replaced by ADD_8288

//KaratsubaCore_473 replaced by KaratsubaCore_1438

//KaratsubaCore_472 replaced by KaratsubaCore_1435

//KaratsubaCore_471 replaced by KaratsubaCore_1438

//BADD_1682 replaced by BADD_2824

//BADD_1681 replaced by BADD_2823

//BADD_1680 replaced by BADD_2822

//ADD_5864 replaced by ADD_11602

//ADD_5863 replaced by ADD_11602

//KaratsubaCore_476 replaced by KaratsubaCore_1437

//KaratsubaCore_475 replaced by KaratsubaCore_1438

//KaratsubaCore_474 replaced by KaratsubaCore_1437

//ADD_5869 replaced by ADD_11595

//ADD_5868 replaced by ADD_11602

//ADD_5867 replaced by ADD_11602

//ADD_5866 replaced by ADD_11602

//ADD_5865 replaced by ADD_11602

//ADD_5874 replaced by ADD_11592

//ADD_5873 replaced by ADD_11602

//ADD_5872 replaced by ADD_11602

//ADD_5871 replaced by ADD_11602

//ADD_5870 replaced by ADD_11602

//ADD_5879 replaced by ADD_11592

//ADD_5878 replaced by ADD_11602

//ADD_5877 replaced by ADD_11602

//ADD_5876 replaced by ADD_11602

//ADD_5875 replaced by ADD_11602

//ADD_5884 replaced by ADD_11595

//ADD_5883 replaced by ADD_11602

//ADD_5882 replaced by ADD_11602

//ADD_5881 replaced by ADD_11602

//ADD_5880 replaced by ADD_11602

//BADD_1686 replaced by BADD_2818

//BADD_1685 replaced by BADD_2820

//BADD_1684 replaced by BADD_2819

//BADD_1683 replaced by BADD_2818

//ADD_5886 replaced by ADD_8288

//ADD_5885 replaced by ADD_8288

//KaratsubaCore_479 replaced by KaratsubaCore_1438

//KaratsubaCore_478 replaced by KaratsubaCore_1435

//KaratsubaCore_477 replaced by KaratsubaCore_1438

//BADD_1690 replaced by BADD_2807

//BADD_1689 replaced by BADD_2809

//BADD_1688 replaced by BADD_2808

//BADD_1687 replaced by BADD_2807

//ADD_5888 replaced by ADD_8267

//ADD_5887 replaced by ADD_8267

//KaratsubaCore_482 replaced by KaratsubaCore_1435

//KaratsubaCore_481 replaced by KaratsubaCore_1426

//KaratsubaCore_480 replaced by KaratsubaCore_1435

//BADD_1694 replaced by BADD_2818

//BADD_1693 replaced by BADD_2820

//BADD_1692 replaced by BADD_2819

//BADD_1691 replaced by BADD_2818

//ADD_5890 replaced by ADD_8288

//ADD_5889 replaced by ADD_8288

//KaratsubaCore_485 replaced by KaratsubaCore_1438

//KaratsubaCore_484 replaced by KaratsubaCore_1435

//KaratsubaCore_483 replaced by KaratsubaCore_1438

//ADD_5896 replaced by ADD_11602

//ADD_5895 replaced by ADD_11602

//ADD_5894 replaced by ADD_11602

//ADD_5893 replaced by ADD_11602

//ADD_5892 replaced by ADD_11602

//ADD_5891 replaced by ADD_11602

//ADD_5901 replaced by ADD_11601

//ADD_5900 replaced by ADD_11602

//ADD_5899 replaced by ADD_11602

//ADD_5898 replaced by ADD_11602

//ADD_5897 replaced by ADD_11602

//ADD_5905 replaced by ADD_11602

//ADD_5904 replaced by ADD_11602

//ADD_5903 replaced by ADD_11602

//ADD_5902 replaced by ADD_11602

//BADD_1697 replaced by BADD_2824

//BADD_1696 replaced by BADD_2823

//BADD_1695 replaced by BADD_2822

//ADD_5907 replaced by ADD_11602

//ADD_5906 replaced by ADD_11602

//KaratsubaCore_488 replaced by KaratsubaCore_1437

//KaratsubaCore_487 replaced by KaratsubaCore_1438

//KaratsubaCore_486 replaced by KaratsubaCore_1437

//BADD_1701 replaced by BADD_2818

//BADD_1700 replaced by BADD_2820

//BADD_1699 replaced by BADD_2819

//BADD_1698 replaced by BADD_2818

//ADD_5909 replaced by ADD_8288

//ADD_5908 replaced by ADD_8288

//KaratsubaCore_491 replaced by KaratsubaCore_1438

//KaratsubaCore_490 replaced by KaratsubaCore_1435

//KaratsubaCore_489 replaced by KaratsubaCore_1438

//BADD_1704 replaced by BADD_2824

//BADD_1703 replaced by BADD_2823

//BADD_1702 replaced by BADD_2822

//ADD_5911 replaced by ADD_11602

//ADD_5910 replaced by ADD_11602

//KaratsubaCore_494 replaced by KaratsubaCore_1437

//KaratsubaCore_493 replaced by KaratsubaCore_1438

//KaratsubaCore_492 replaced by KaratsubaCore_1437

//ADD_5917 replaced by ADD_11602

//ADD_5916 replaced by ADD_11602

//ADD_5915 replaced by ADD_11602

//ADD_5914 replaced by ADD_11602

//ADD_5913 replaced by ADD_11602

//ADD_5912 replaced by ADD_11602

//ADD_5922 replaced by ADD_11601

//ADD_5921 replaced by ADD_11602

//ADD_5920 replaced by ADD_11602

//ADD_5919 replaced by ADD_11602

//ADD_5918 replaced by ADD_11602

//ADD_5926 replaced by ADD_11602

//ADD_5925 replaced by ADD_11602

//ADD_5924 replaced by ADD_11602

//ADD_5923 replaced by ADD_11602

//BADD_1707 replaced by BADD_2824

//BADD_1706 replaced by BADD_2823

//BADD_1705 replaced by BADD_2822

//ADD_5928 replaced by ADD_11602

//ADD_5927 replaced by ADD_11602

//KaratsubaCore_497 replaced by KaratsubaCore_1437

//KaratsubaCore_496 replaced by KaratsubaCore_1438

//KaratsubaCore_495 replaced by KaratsubaCore_1437

//BADD_1711 replaced by BADD_2818

//BADD_1710 replaced by BADD_2820

//BADD_1709 replaced by BADD_2819

//BADD_1708 replaced by BADD_2818

//ADD_5930 replaced by ADD_8288

//ADD_5929 replaced by ADD_8288

//KaratsubaCore_500 replaced by KaratsubaCore_1438

//KaratsubaCore_499 replaced by KaratsubaCore_1435

//KaratsubaCore_498 replaced by KaratsubaCore_1438

//BADD_1714 replaced by BADD_2824

//BADD_1713 replaced by BADD_2823

//BADD_1712 replaced by BADD_2822

//ADD_5932 replaced by ADD_11602

//ADD_5931 replaced by ADD_11602

//KaratsubaCore_503 replaced by KaratsubaCore_1437

//KaratsubaCore_502 replaced by KaratsubaCore_1438

//KaratsubaCore_501 replaced by KaratsubaCore_1437

//ADD_5937 replaced by ADD_11595

//ADD_5936 replaced by ADD_11602

//ADD_5935 replaced by ADD_11602

//ADD_5934 replaced by ADD_11602

//ADD_5933 replaced by ADD_11602

//ADD_5942 replaced by ADD_11592

//ADD_5941 replaced by ADD_11602

//ADD_5940 replaced by ADD_11602

//ADD_5939 replaced by ADD_11602

//ADD_5938 replaced by ADD_11602

//ADD_5947 replaced by ADD_11592

//ADD_5946 replaced by ADD_11602

//ADD_5945 replaced by ADD_11602

//ADD_5944 replaced by ADD_11602

//ADD_5943 replaced by ADD_11602

//ADD_5952 replaced by ADD_11595

//ADD_5951 replaced by ADD_11602

//ADD_5950 replaced by ADD_11602

//ADD_5949 replaced by ADD_11602

//ADD_5948 replaced by ADD_11602

//BADD_1718 replaced by BADD_2818

//BADD_1717 replaced by BADD_2820

//BADD_1716 replaced by BADD_2819

//BADD_1715 replaced by BADD_2818

//ADD_5954 replaced by ADD_8288

//ADD_5953 replaced by ADD_8288

//KaratsubaCore_506 replaced by KaratsubaCore_1438

//KaratsubaCore_505 replaced by KaratsubaCore_1435

//KaratsubaCore_504 replaced by KaratsubaCore_1438

//BADD_1722 replaced by BADD_2807

//BADD_1721 replaced by BADD_2809

//BADD_1720 replaced by BADD_2808

//BADD_1719 replaced by BADD_2807

//ADD_5956 replaced by ADD_8267

//ADD_5955 replaced by ADD_8267

//KaratsubaCore_509 replaced by KaratsubaCore_1435

//KaratsubaCore_508 replaced by KaratsubaCore_1426

//KaratsubaCore_507 replaced by KaratsubaCore_1435

//BADD_1726 replaced by BADD_2818

//BADD_1725 replaced by BADD_2820

//BADD_1724 replaced by BADD_2819

//BADD_1723 replaced by BADD_2818

//ADD_5958 replaced by ADD_8288

//ADD_5957 replaced by ADD_8288

//KaratsubaCore_512 replaced by KaratsubaCore_1438

//KaratsubaCore_511 replaced by KaratsubaCore_1435

//KaratsubaCore_510 replaced by KaratsubaCore_1438

//ADD_5964 replaced by ADD_11602

//ADD_5963 replaced by ADD_11602

//ADD_5962 replaced by ADD_11602

//ADD_5961 replaced by ADD_11602

//ADD_5960 replaced by ADD_11602

//ADD_5959 replaced by ADD_11602

//ADD_5969 replaced by ADD_11601

//ADD_5968 replaced by ADD_11602

//ADD_5967 replaced by ADD_11602

//ADD_5966 replaced by ADD_11602

//ADD_5965 replaced by ADD_11602

//ADD_5973 replaced by ADD_11602

//ADD_5972 replaced by ADD_11602

//ADD_5971 replaced by ADD_11602

//ADD_5970 replaced by ADD_11602

//BADD_1729 replaced by BADD_2824

//BADD_1728 replaced by BADD_2823

//BADD_1727 replaced by BADD_2822

//ADD_5975 replaced by ADD_11602

//ADD_5974 replaced by ADD_11602

//KaratsubaCore_515 replaced by KaratsubaCore_1437

//KaratsubaCore_514 replaced by KaratsubaCore_1438

//KaratsubaCore_513 replaced by KaratsubaCore_1437

//BADD_1733 replaced by BADD_2818

//BADD_1732 replaced by BADD_2820

//BADD_1731 replaced by BADD_2819

//BADD_1730 replaced by BADD_2818

//ADD_5977 replaced by ADD_8288

//ADD_5976 replaced by ADD_8288

//KaratsubaCore_518 replaced by KaratsubaCore_1438

//KaratsubaCore_517 replaced by KaratsubaCore_1435

//KaratsubaCore_516 replaced by KaratsubaCore_1438

//BADD_1736 replaced by BADD_2824

//BADD_1735 replaced by BADD_2823

//BADD_1734 replaced by BADD_2822

//ADD_5979 replaced by ADD_11602

//ADD_5978 replaced by ADD_11602

//KaratsubaCore_521 replaced by KaratsubaCore_1437

//KaratsubaCore_520 replaced by KaratsubaCore_1438

//KaratsubaCore_519 replaced by KaratsubaCore_1437

//ADD_5985 replaced by ADD_11602

//ADD_5984 replaced by ADD_11602

//ADD_5983 replaced by ADD_11602

//ADD_5982 replaced by ADD_11602

//ADD_5981 replaced by ADD_11602

//ADD_5980 replaced by ADD_11602

//ADD_5990 replaced by ADD_11601

//ADD_5989 replaced by ADD_11602

//ADD_5988 replaced by ADD_11602

//ADD_5987 replaced by ADD_11602

//ADD_5986 replaced by ADD_11602

//ADD_5994 replaced by ADD_11602

//ADD_5993 replaced by ADD_11602

//ADD_5992 replaced by ADD_11602

//ADD_5991 replaced by ADD_11602

//BADD_1739 replaced by BADD_2824

//BADD_1738 replaced by BADD_2823

//BADD_1737 replaced by BADD_2822

//ADD_5996 replaced by ADD_11602

//ADD_5995 replaced by ADD_11602

//KaratsubaCore_524 replaced by KaratsubaCore_1437

//KaratsubaCore_523 replaced by KaratsubaCore_1438

//KaratsubaCore_522 replaced by KaratsubaCore_1437

//BADD_1743 replaced by BADD_2818

//BADD_1742 replaced by BADD_2820

//BADD_1741 replaced by BADD_2819

//BADD_1740 replaced by BADD_2818

//ADD_5998 replaced by ADD_8288

//ADD_5997 replaced by ADD_8288

//KaratsubaCore_527 replaced by KaratsubaCore_1438

//KaratsubaCore_526 replaced by KaratsubaCore_1435

//KaratsubaCore_525 replaced by KaratsubaCore_1438

//BADD_1746 replaced by BADD_2824

//BADD_1745 replaced by BADD_2823

//BADD_1744 replaced by BADD_2822

//ADD_6000 replaced by ADD_11602

//ADD_5999 replaced by ADD_11602

//KaratsubaCore_530 replaced by KaratsubaCore_1437

//KaratsubaCore_529 replaced by KaratsubaCore_1438

//KaratsubaCore_528 replaced by KaratsubaCore_1437

//ADD_6005 replaced by ADD_11595

//ADD_6004 replaced by ADD_11602

//ADD_6003 replaced by ADD_11602

//ADD_6002 replaced by ADD_11602

//ADD_6001 replaced by ADD_11602

//ADD_6010 replaced by ADD_11592

//ADD_6009 replaced by ADD_11602

//ADD_6008 replaced by ADD_11602

//ADD_6007 replaced by ADD_11602

//ADD_6006 replaced by ADD_11602

//ADD_6015 replaced by ADD_11592

//ADD_6014 replaced by ADD_11602

//ADD_6013 replaced by ADD_11602

//ADD_6012 replaced by ADD_11602

//ADD_6011 replaced by ADD_11602

//ADD_6020 replaced by ADD_11595

//ADD_6019 replaced by ADD_11602

//ADD_6018 replaced by ADD_11602

//ADD_6017 replaced by ADD_11602

//ADD_6016 replaced by ADD_11602

//BADD_1750 replaced by BADD_2818

//BADD_1749 replaced by BADD_2820

//BADD_1748 replaced by BADD_2819

//BADD_1747 replaced by BADD_2818

//ADD_6022 replaced by ADD_8288

//ADD_6021 replaced by ADD_8288

//KaratsubaCore_533 replaced by KaratsubaCore_1438

//KaratsubaCore_532 replaced by KaratsubaCore_1435

//KaratsubaCore_531 replaced by KaratsubaCore_1438

//BADD_1754 replaced by BADD_2807

//BADD_1753 replaced by BADD_2809

//BADD_1752 replaced by BADD_2808

//BADD_1751 replaced by BADD_2807

//ADD_6024 replaced by ADD_8267

//ADD_6023 replaced by ADD_8267

//KaratsubaCore_536 replaced by KaratsubaCore_1435

//KaratsubaCore_535 replaced by KaratsubaCore_1426

//KaratsubaCore_534 replaced by KaratsubaCore_1435

//BADD_1758 replaced by BADD_2818

//BADD_1757 replaced by BADD_2820

//BADD_1756 replaced by BADD_2819

//BADD_1755 replaced by BADD_2818

//ADD_6026 replaced by ADD_8288

//ADD_6025 replaced by ADD_8288

//KaratsubaCore_539 replaced by KaratsubaCore_1438

//KaratsubaCore_538 replaced by KaratsubaCore_1435

//KaratsubaCore_537 replaced by KaratsubaCore_1438

//ADD_6032 replaced by ADD_11602

//ADD_6031 replaced by ADD_11602

//ADD_6030 replaced by ADD_11602

//ADD_6029 replaced by ADD_11602

//ADD_6028 replaced by ADD_11602

//ADD_6027 replaced by ADD_11602

//ADD_6037 replaced by ADD_11601

//ADD_6036 replaced by ADD_11602

//ADD_6035 replaced by ADD_11602

//ADD_6034 replaced by ADD_11602

//ADD_6033 replaced by ADD_11602

//ADD_6041 replaced by ADD_11602

//ADD_6040 replaced by ADD_11602

//ADD_6039 replaced by ADD_11602

//ADD_6038 replaced by ADD_11602

//BADD_1761 replaced by BADD_2824

//BADD_1760 replaced by BADD_2823

//BADD_1759 replaced by BADD_2822

//ADD_6043 replaced by ADD_11602

//ADD_6042 replaced by ADD_11602

//KaratsubaCore_542 replaced by KaratsubaCore_1437

//KaratsubaCore_541 replaced by KaratsubaCore_1438

//KaratsubaCore_540 replaced by KaratsubaCore_1437

//BADD_1765 replaced by BADD_2818

//BADD_1764 replaced by BADD_2820

//BADD_1763 replaced by BADD_2819

//BADD_1762 replaced by BADD_2818

//ADD_6045 replaced by ADD_8288

//ADD_6044 replaced by ADD_8288

//KaratsubaCore_545 replaced by KaratsubaCore_1438

//KaratsubaCore_544 replaced by KaratsubaCore_1435

//KaratsubaCore_543 replaced by KaratsubaCore_1438

//BADD_1768 replaced by BADD_2824

//BADD_1767 replaced by BADD_2823

//BADD_1766 replaced by BADD_2822

//ADD_6047 replaced by ADD_11602

//ADD_6046 replaced by ADD_11602

//KaratsubaCore_548 replaced by KaratsubaCore_1437

//KaratsubaCore_547 replaced by KaratsubaCore_1438

//KaratsubaCore_546 replaced by KaratsubaCore_1437

//ADD_6053 replaced by ADD_11602

//ADD_6052 replaced by ADD_11602

//ADD_6051 replaced by ADD_11602

//ADD_6050 replaced by ADD_11602

//ADD_6049 replaced by ADD_11602

//ADD_6048 replaced by ADD_11602

//ADD_6058 replaced by ADD_11601

//ADD_6057 replaced by ADD_11602

//ADD_6056 replaced by ADD_11602

//ADD_6055 replaced by ADD_11602

//ADD_6054 replaced by ADD_11602

//ADD_6062 replaced by ADD_11602

//ADD_6061 replaced by ADD_11602

//ADD_6060 replaced by ADD_11602

//ADD_6059 replaced by ADD_11602

//BADD_1771 replaced by BADD_2824

//BADD_1770 replaced by BADD_2823

//BADD_1769 replaced by BADD_2822

//ADD_6064 replaced by ADD_11602

//ADD_6063 replaced by ADD_11602

//KaratsubaCore_551 replaced by KaratsubaCore_1437

//KaratsubaCore_550 replaced by KaratsubaCore_1438

//KaratsubaCore_549 replaced by KaratsubaCore_1437

//BADD_1775 replaced by BADD_2818

//BADD_1774 replaced by BADD_2820

//BADD_1773 replaced by BADD_2819

//BADD_1772 replaced by BADD_2818

//ADD_6066 replaced by ADD_8288

//ADD_6065 replaced by ADD_8288

//KaratsubaCore_554 replaced by KaratsubaCore_1438

//KaratsubaCore_553 replaced by KaratsubaCore_1435

//KaratsubaCore_552 replaced by KaratsubaCore_1438

//BADD_1778 replaced by BADD_2824

//BADD_1777 replaced by BADD_2823

//BADD_1776 replaced by BADD_2822

//ADD_6068 replaced by ADD_11602

//ADD_6067 replaced by ADD_11602

//KaratsubaCore_557 replaced by KaratsubaCore_1437

//KaratsubaCore_556 replaced by KaratsubaCore_1438

//KaratsubaCore_555 replaced by KaratsubaCore_1437

//ADD_6073 replaced by ADD_11595

//ADD_6072 replaced by ADD_11602

//ADD_6071 replaced by ADD_11602

//ADD_6070 replaced by ADD_11602

//ADD_6069 replaced by ADD_11602

//ADD_6078 replaced by ADD_11592

//ADD_6077 replaced by ADD_11602

//ADD_6076 replaced by ADD_11602

//ADD_6075 replaced by ADD_11602

//ADD_6074 replaced by ADD_11602

//ADD_6083 replaced by ADD_11592

//ADD_6082 replaced by ADD_11602

//ADD_6081 replaced by ADD_11602

//ADD_6080 replaced by ADD_11602

//ADD_6079 replaced by ADD_11602

//ADD_6088 replaced by ADD_11595

//ADD_6087 replaced by ADD_11602

//ADD_6086 replaced by ADD_11602

//ADD_6085 replaced by ADD_11602

//ADD_6084 replaced by ADD_11602

//BADD_1782 replaced by BADD_2818

//BADD_1781 replaced by BADD_2820

//BADD_1780 replaced by BADD_2819

//BADD_1779 replaced by BADD_2818

//ADD_6090 replaced by ADD_8288

//ADD_6089 replaced by ADD_8288

//KaratsubaCore_560 replaced by KaratsubaCore_1438

//KaratsubaCore_559 replaced by KaratsubaCore_1435

//KaratsubaCore_558 replaced by KaratsubaCore_1438

//BADD_1786 replaced by BADD_2807

//BADD_1785 replaced by BADD_2809

//BADD_1784 replaced by BADD_2808

//BADD_1783 replaced by BADD_2807

//ADD_6092 replaced by ADD_8267

//ADD_6091 replaced by ADD_8267

//KaratsubaCore_563 replaced by KaratsubaCore_1435

//KaratsubaCore_562 replaced by KaratsubaCore_1426

//KaratsubaCore_561 replaced by KaratsubaCore_1435

//BADD_1790 replaced by BADD_2818

//BADD_1789 replaced by BADD_2820

//BADD_1788 replaced by BADD_2819

//BADD_1787 replaced by BADD_2818

//ADD_6094 replaced by ADD_8288

//ADD_6093 replaced by ADD_8288

//KaratsubaCore_566 replaced by KaratsubaCore_1438

//KaratsubaCore_565 replaced by KaratsubaCore_1435

//KaratsubaCore_564 replaced by KaratsubaCore_1438

//ADD_6100 replaced by ADD_11602

//ADD_6099 replaced by ADD_11602

//ADD_6098 replaced by ADD_11602

//ADD_6097 replaced by ADD_11602

//ADD_6096 replaced by ADD_11602

//ADD_6095 replaced by ADD_11602

//ADD_6105 replaced by ADD_11601

//ADD_6104 replaced by ADD_11602

//ADD_6103 replaced by ADD_11602

//ADD_6102 replaced by ADD_11602

//ADD_6101 replaced by ADD_11602

//ADD_6109 replaced by ADD_11602

//ADD_6108 replaced by ADD_11602

//ADD_6107 replaced by ADD_11602

//ADD_6106 replaced by ADD_11602

//BADD_1793 replaced by BADD_2824

//BADD_1792 replaced by BADD_2823

//BADD_1791 replaced by BADD_2822

//ADD_6111 replaced by ADD_11602

//ADD_6110 replaced by ADD_11602

//KaratsubaCore_569 replaced by KaratsubaCore_1437

//KaratsubaCore_568 replaced by KaratsubaCore_1438

//KaratsubaCore_567 replaced by KaratsubaCore_1437

//BADD_1797 replaced by BADD_2818

//BADD_1796 replaced by BADD_2820

//BADD_1795 replaced by BADD_2819

//BADD_1794 replaced by BADD_2818

//ADD_6113 replaced by ADD_8288

//ADD_6112 replaced by ADD_8288

//KaratsubaCore_572 replaced by KaratsubaCore_1438

//KaratsubaCore_571 replaced by KaratsubaCore_1435

//KaratsubaCore_570 replaced by KaratsubaCore_1438

//BADD_1800 replaced by BADD_2824

//BADD_1799 replaced by BADD_2823

//BADD_1798 replaced by BADD_2822

//ADD_6115 replaced by ADD_11602

//ADD_6114 replaced by ADD_11602

//KaratsubaCore_575 replaced by KaratsubaCore_1437

//KaratsubaCore_574 replaced by KaratsubaCore_1438

//KaratsubaCore_573 replaced by KaratsubaCore_1437

//ADD_6121 replaced by ADD_11602

//ADD_6120 replaced by ADD_11602

//ADD_6119 replaced by ADD_11602

//ADD_6118 replaced by ADD_11602

//ADD_6117 replaced by ADD_11602

//ADD_6116 replaced by ADD_11602

//ADD_6126 replaced by ADD_11601

//ADD_6125 replaced by ADD_11602

//ADD_6124 replaced by ADD_11602

//ADD_6123 replaced by ADD_11602

//ADD_6122 replaced by ADD_11602

//ADD_6130 replaced by ADD_11602

//ADD_6129 replaced by ADD_11602

//ADD_6128 replaced by ADD_11602

//ADD_6127 replaced by ADD_11602

//BADD_1803 replaced by BADD_2824

//BADD_1802 replaced by BADD_2823

//BADD_1801 replaced by BADD_2822

//ADD_6132 replaced by ADD_11602

//ADD_6131 replaced by ADD_11602

//KaratsubaCore_578 replaced by KaratsubaCore_1437

//KaratsubaCore_577 replaced by KaratsubaCore_1438

//KaratsubaCore_576 replaced by KaratsubaCore_1437

//BADD_1807 replaced by BADD_2818

//BADD_1806 replaced by BADD_2820

//BADD_1805 replaced by BADD_2819

//BADD_1804 replaced by BADD_2818

//ADD_6134 replaced by ADD_8288

//ADD_6133 replaced by ADD_8288

//KaratsubaCore_581 replaced by KaratsubaCore_1438

//KaratsubaCore_580 replaced by KaratsubaCore_1435

//KaratsubaCore_579 replaced by KaratsubaCore_1438

//BADD_1810 replaced by BADD_2824

//BADD_1809 replaced by BADD_2823

//BADD_1808 replaced by BADD_2822

//ADD_6136 replaced by ADD_11602

//ADD_6135 replaced by ADD_11602

//KaratsubaCore_584 replaced by KaratsubaCore_1437

//KaratsubaCore_583 replaced by KaratsubaCore_1438

//KaratsubaCore_582 replaced by KaratsubaCore_1437

//ADD_6141 replaced by ADD_11595

//ADD_6140 replaced by ADD_11602

//ADD_6139 replaced by ADD_11602

//ADD_6138 replaced by ADD_11602

//ADD_6137 replaced by ADD_11602

//ADD_6146 replaced by ADD_11592

//ADD_6145 replaced by ADD_11602

//ADD_6144 replaced by ADD_11602

//ADD_6143 replaced by ADD_11602

//ADD_6142 replaced by ADD_11602

//ADD_6151 replaced by ADD_11592

//ADD_6150 replaced by ADD_11602

//ADD_6149 replaced by ADD_11602

//ADD_6148 replaced by ADD_11602

//ADD_6147 replaced by ADD_11602

//ADD_6156 replaced by ADD_11595

//ADD_6155 replaced by ADD_11602

//ADD_6154 replaced by ADD_11602

//ADD_6153 replaced by ADD_11602

//ADD_6152 replaced by ADD_11602

//BADD_1814 replaced by BADD_2818

//BADD_1813 replaced by BADD_2820

//BADD_1812 replaced by BADD_2819

//BADD_1811 replaced by BADD_2818

//ADD_6158 replaced by ADD_8288

//ADD_6157 replaced by ADD_8288

//KaratsubaCore_587 replaced by KaratsubaCore_1438

//KaratsubaCore_586 replaced by KaratsubaCore_1435

//KaratsubaCore_585 replaced by KaratsubaCore_1438

//BADD_1818 replaced by BADD_2807

//BADD_1817 replaced by BADD_2809

//BADD_1816 replaced by BADD_2808

//BADD_1815 replaced by BADD_2807

//ADD_6160 replaced by ADD_8267

//ADD_6159 replaced by ADD_8267

//KaratsubaCore_590 replaced by KaratsubaCore_1435

//KaratsubaCore_589 replaced by KaratsubaCore_1426

//KaratsubaCore_588 replaced by KaratsubaCore_1435

//BADD_1822 replaced by BADD_2818

//BADD_1821 replaced by BADD_2820

//BADD_1820 replaced by BADD_2819

//BADD_1819 replaced by BADD_2818

//ADD_6162 replaced by ADD_8288

//ADD_6161 replaced by ADD_8288

//KaratsubaCore_593 replaced by KaratsubaCore_1438

//KaratsubaCore_592 replaced by KaratsubaCore_1435

//KaratsubaCore_591 replaced by KaratsubaCore_1438

//ADD_6168 replaced by ADD_11602

//ADD_6167 replaced by ADD_11602

//ADD_6166 replaced by ADD_11602

//ADD_6165 replaced by ADD_11602

//ADD_6164 replaced by ADD_11602

//ADD_6163 replaced by ADD_11602

//ADD_6173 replaced by ADD_11601

//ADD_6172 replaced by ADD_11602

//ADD_6171 replaced by ADD_11602

//ADD_6170 replaced by ADD_11602

//ADD_6169 replaced by ADD_11602

//ADD_6177 replaced by ADD_11602

//ADD_6176 replaced by ADD_11602

//ADD_6175 replaced by ADD_11602

//ADD_6174 replaced by ADD_11602

//BADD_1825 replaced by BADD_2824

//BADD_1824 replaced by BADD_2823

//BADD_1823 replaced by BADD_2822

//ADD_6179 replaced by ADD_11602

//ADD_6178 replaced by ADD_11602

//KaratsubaCore_596 replaced by KaratsubaCore_1437

//KaratsubaCore_595 replaced by KaratsubaCore_1438

//KaratsubaCore_594 replaced by KaratsubaCore_1437

//BADD_1829 replaced by BADD_2818

//BADD_1828 replaced by BADD_2820

//BADD_1827 replaced by BADD_2819

//BADD_1826 replaced by BADD_2818

//ADD_6181 replaced by ADD_8288

//ADD_6180 replaced by ADD_8288

//KaratsubaCore_599 replaced by KaratsubaCore_1438

//KaratsubaCore_598 replaced by KaratsubaCore_1435

//KaratsubaCore_597 replaced by KaratsubaCore_1438

//BADD_1832 replaced by BADD_2824

//BADD_1831 replaced by BADD_2823

//BADD_1830 replaced by BADD_2822

//ADD_6183 replaced by ADD_11602

//ADD_6182 replaced by ADD_11602

//KaratsubaCore_602 replaced by KaratsubaCore_1437

//KaratsubaCore_601 replaced by KaratsubaCore_1438

//KaratsubaCore_600 replaced by KaratsubaCore_1437

//ADD_6189 replaced by ADD_11602

//ADD_6188 replaced by ADD_11602

//ADD_6187 replaced by ADD_11602

//ADD_6186 replaced by ADD_11602

//ADD_6185 replaced by ADD_11602

//ADD_6184 replaced by ADD_11602

//ADD_6194 replaced by ADD_11601

//ADD_6193 replaced by ADD_11602

//ADD_6192 replaced by ADD_11602

//ADD_6191 replaced by ADD_11602

//ADD_6190 replaced by ADD_11602

//ADD_6198 replaced by ADD_11602

//ADD_6197 replaced by ADD_11602

//ADD_6196 replaced by ADD_11602

//ADD_6195 replaced by ADD_11602

//BADD_1835 replaced by BADD_2824

//BADD_1834 replaced by BADD_2823

//BADD_1833 replaced by BADD_2822

//ADD_6200 replaced by ADD_11602

//ADD_6199 replaced by ADD_11602

//KaratsubaCore_605 replaced by KaratsubaCore_1437

//KaratsubaCore_604 replaced by KaratsubaCore_1438

//KaratsubaCore_603 replaced by KaratsubaCore_1437

//BADD_1839 replaced by BADD_2818

//BADD_1838 replaced by BADD_2820

//BADD_1837 replaced by BADD_2819

//BADD_1836 replaced by BADD_2818

//ADD_6202 replaced by ADD_8288

//ADD_6201 replaced by ADD_8288

//KaratsubaCore_608 replaced by KaratsubaCore_1438

//KaratsubaCore_607 replaced by KaratsubaCore_1435

//KaratsubaCore_606 replaced by KaratsubaCore_1438

//BADD_1842 replaced by BADD_2824

//BADD_1841 replaced by BADD_2823

//BADD_1840 replaced by BADD_2822

//ADD_6204 replaced by ADD_11602

//ADD_6203 replaced by ADD_11602

//KaratsubaCore_611 replaced by KaratsubaCore_1437

//KaratsubaCore_610 replaced by KaratsubaCore_1438

//KaratsubaCore_609 replaced by KaratsubaCore_1437

//ADD_6209 replaced by ADD_11595

//ADD_6208 replaced by ADD_11602

//ADD_6207 replaced by ADD_11602

//ADD_6206 replaced by ADD_11602

//ADD_6205 replaced by ADD_11602

//ADD_6214 replaced by ADD_11592

//ADD_6213 replaced by ADD_11602

//ADD_6212 replaced by ADD_11602

//ADD_6211 replaced by ADD_11602

//ADD_6210 replaced by ADD_11602

//ADD_6219 replaced by ADD_11592

//ADD_6218 replaced by ADD_11602

//ADD_6217 replaced by ADD_11602

//ADD_6216 replaced by ADD_11602

//ADD_6215 replaced by ADD_11602

//ADD_6224 replaced by ADD_11595

//ADD_6223 replaced by ADD_11602

//ADD_6222 replaced by ADD_11602

//ADD_6221 replaced by ADD_11602

//ADD_6220 replaced by ADD_11602

//BADD_1846 replaced by BADD_2818

//BADD_1845 replaced by BADD_2820

//BADD_1844 replaced by BADD_2819

//BADD_1843 replaced by BADD_2818

//ADD_6226 replaced by ADD_8288

//ADD_6225 replaced by ADD_8288

//KaratsubaCore_614 replaced by KaratsubaCore_1438

//KaratsubaCore_613 replaced by KaratsubaCore_1435

//KaratsubaCore_612 replaced by KaratsubaCore_1438

//BADD_1850 replaced by BADD_2807

//BADD_1849 replaced by BADD_2809

//BADD_1848 replaced by BADD_2808

//BADD_1847 replaced by BADD_2807

//ADD_6228 replaced by ADD_8267

//ADD_6227 replaced by ADD_8267

//KaratsubaCore_617 replaced by KaratsubaCore_1435

//KaratsubaCore_616 replaced by KaratsubaCore_1426

//KaratsubaCore_615 replaced by KaratsubaCore_1435

//BADD_1854 replaced by BADD_2818

//BADD_1853 replaced by BADD_2820

//BADD_1852 replaced by BADD_2819

//BADD_1851 replaced by BADD_2818

//ADD_6230 replaced by ADD_8288

//ADD_6229 replaced by ADD_8288

//KaratsubaCore_620 replaced by KaratsubaCore_1438

//KaratsubaCore_619 replaced by KaratsubaCore_1435

//KaratsubaCore_618 replaced by KaratsubaCore_1438

//ADD_6236 replaced by ADD_11602

//ADD_6235 replaced by ADD_11602

//ADD_6234 replaced by ADD_11602

//ADD_6233 replaced by ADD_11602

//ADD_6232 replaced by ADD_11602

//ADD_6231 replaced by ADD_11602

//ADD_6241 replaced by ADD_11601

//ADD_6240 replaced by ADD_11602

//ADD_6239 replaced by ADD_11602

//ADD_6238 replaced by ADD_11602

//ADD_6237 replaced by ADD_11602

//ADD_6245 replaced by ADD_11602

//ADD_6244 replaced by ADD_11602

//ADD_6243 replaced by ADD_11602

//ADD_6242 replaced by ADD_11602

//BADD_1857 replaced by BADD_2824

//BADD_1856 replaced by BADD_2823

//BADD_1855 replaced by BADD_2822

//ADD_6247 replaced by ADD_11602

//ADD_6246 replaced by ADD_11602

//KaratsubaCore_623 replaced by KaratsubaCore_1437

//KaratsubaCore_622 replaced by KaratsubaCore_1438

//KaratsubaCore_621 replaced by KaratsubaCore_1437

//BADD_1861 replaced by BADD_2818

//BADD_1860 replaced by BADD_2820

//BADD_1859 replaced by BADD_2819

//BADD_1858 replaced by BADD_2818

//ADD_6249 replaced by ADD_8288

//ADD_6248 replaced by ADD_8288

//KaratsubaCore_626 replaced by KaratsubaCore_1438

//KaratsubaCore_625 replaced by KaratsubaCore_1435

//KaratsubaCore_624 replaced by KaratsubaCore_1438

//BADD_1864 replaced by BADD_2824

//BADD_1863 replaced by BADD_2823

//BADD_1862 replaced by BADD_2822

//ADD_6251 replaced by ADD_11602

//ADD_6250 replaced by ADD_11602

//KaratsubaCore_629 replaced by KaratsubaCore_1437

//KaratsubaCore_628 replaced by KaratsubaCore_1438

//KaratsubaCore_627 replaced by KaratsubaCore_1437

//ADD_6257 replaced by ADD_11602

//ADD_6256 replaced by ADD_11602

//ADD_6255 replaced by ADD_11602

//ADD_6254 replaced by ADD_11602

//ADD_6253 replaced by ADD_11602

//ADD_6252 replaced by ADD_11602

//ADD_6262 replaced by ADD_11601

//ADD_6261 replaced by ADD_11602

//ADD_6260 replaced by ADD_11602

//ADD_6259 replaced by ADD_11602

//ADD_6258 replaced by ADD_11602

//ADD_6266 replaced by ADD_11602

//ADD_6265 replaced by ADD_11602

//ADD_6264 replaced by ADD_11602

//ADD_6263 replaced by ADD_11602

//BADD_1867 replaced by BADD_2824

//BADD_1866 replaced by BADD_2823

//BADD_1865 replaced by BADD_2822

//ADD_6268 replaced by ADD_11602

//ADD_6267 replaced by ADD_11602

//KaratsubaCore_632 replaced by KaratsubaCore_1437

//KaratsubaCore_631 replaced by KaratsubaCore_1438

//KaratsubaCore_630 replaced by KaratsubaCore_1437

//BADD_1871 replaced by BADD_2818

//BADD_1870 replaced by BADD_2820

//BADD_1869 replaced by BADD_2819

//BADD_1868 replaced by BADD_2818

//ADD_6270 replaced by ADD_8288

//ADD_6269 replaced by ADD_8288

//KaratsubaCore_635 replaced by KaratsubaCore_1438

//KaratsubaCore_634 replaced by KaratsubaCore_1435

//KaratsubaCore_633 replaced by KaratsubaCore_1438

//BADD_1874 replaced by BADD_2824

//BADD_1873 replaced by BADD_2823

//BADD_1872 replaced by BADD_2822

//ADD_6272 replaced by ADD_11602

//ADD_6271 replaced by ADD_11602

//KaratsubaCore_638 replaced by KaratsubaCore_1437

//KaratsubaCore_637 replaced by KaratsubaCore_1438

//KaratsubaCore_636 replaced by KaratsubaCore_1437

//ADD_6277 replaced by ADD_11595

//ADD_6276 replaced by ADD_11602

//ADD_6275 replaced by ADD_11602

//ADD_6274 replaced by ADD_11602

//ADD_6273 replaced by ADD_11602

//ADD_6282 replaced by ADD_11592

//ADD_6281 replaced by ADD_11602

//ADD_6280 replaced by ADD_11602

//ADD_6279 replaced by ADD_11602

//ADD_6278 replaced by ADD_11602

//ADD_6287 replaced by ADD_11592

//ADD_6286 replaced by ADD_11602

//ADD_6285 replaced by ADD_11602

//ADD_6284 replaced by ADD_11602

//ADD_6283 replaced by ADD_11602

//ADD_6292 replaced by ADD_11595

//ADD_6291 replaced by ADD_11602

//ADD_6290 replaced by ADD_11602

//ADD_6289 replaced by ADD_11602

//ADD_6288 replaced by ADD_11602

//BADD_1878 replaced by BADD_2818

//BADD_1877 replaced by BADD_2820

//BADD_1876 replaced by BADD_2819

//BADD_1875 replaced by BADD_2818

//ADD_6294 replaced by ADD_8288

//ADD_6293 replaced by ADD_8288

//KaratsubaCore_641 replaced by KaratsubaCore_1438

//KaratsubaCore_640 replaced by KaratsubaCore_1435

//KaratsubaCore_639 replaced by KaratsubaCore_1438

//BADD_1882 replaced by BADD_2807

//BADD_1881 replaced by BADD_2809

//BADD_1880 replaced by BADD_2808

//BADD_1879 replaced by BADD_2807

//ADD_6296 replaced by ADD_8267

//ADD_6295 replaced by ADD_8267

//KaratsubaCore_644 replaced by KaratsubaCore_1435

//KaratsubaCore_643 replaced by KaratsubaCore_1426

//KaratsubaCore_642 replaced by KaratsubaCore_1435

//BADD_1886 replaced by BADD_2818

//BADD_1885 replaced by BADD_2820

//BADD_1884 replaced by BADD_2819

//BADD_1883 replaced by BADD_2818

//ADD_6298 replaced by ADD_8288

//ADD_6297 replaced by ADD_8288

//KaratsubaCore_647 replaced by KaratsubaCore_1438

//KaratsubaCore_646 replaced by KaratsubaCore_1435

//KaratsubaCore_645 replaced by KaratsubaCore_1438

//ADD_6304 replaced by ADD_11602

//ADD_6303 replaced by ADD_11602

//ADD_6302 replaced by ADD_11602

//ADD_6301 replaced by ADD_11602

//ADD_6300 replaced by ADD_11602

//ADD_6299 replaced by ADD_11602

//ADD_6309 replaced by ADD_11601

//ADD_6308 replaced by ADD_11602

//ADD_6307 replaced by ADD_11602

//ADD_6306 replaced by ADD_11602

//ADD_6305 replaced by ADD_11602

//ADD_6313 replaced by ADD_11602

//ADD_6312 replaced by ADD_11602

//ADD_6311 replaced by ADD_11602

//ADD_6310 replaced by ADD_11602

//BADD_1889 replaced by BADD_2824

//BADD_1888 replaced by BADD_2823

//BADD_1887 replaced by BADD_2822

//ADD_6315 replaced by ADD_11602

//ADD_6314 replaced by ADD_11602

//KaratsubaCore_650 replaced by KaratsubaCore_1437

//KaratsubaCore_649 replaced by KaratsubaCore_1438

//KaratsubaCore_648 replaced by KaratsubaCore_1437

//BADD_1893 replaced by BADD_2818

//BADD_1892 replaced by BADD_2820

//BADD_1891 replaced by BADD_2819

//BADD_1890 replaced by BADD_2818

//ADD_6317 replaced by ADD_8288

//ADD_6316 replaced by ADD_8288

//KaratsubaCore_653 replaced by KaratsubaCore_1438

//KaratsubaCore_652 replaced by KaratsubaCore_1435

//KaratsubaCore_651 replaced by KaratsubaCore_1438

//BADD_1896 replaced by BADD_2824

//BADD_1895 replaced by BADD_2823

//BADD_1894 replaced by BADD_2822

//ADD_6319 replaced by ADD_11602

//ADD_6318 replaced by ADD_11602

//KaratsubaCore_656 replaced by KaratsubaCore_1437

//KaratsubaCore_655 replaced by KaratsubaCore_1438

//KaratsubaCore_654 replaced by KaratsubaCore_1437

//ADD_6325 replaced by ADD_11602

//ADD_6324 replaced by ADD_11602

//ADD_6323 replaced by ADD_11602

//ADD_6322 replaced by ADD_11602

//ADD_6321 replaced by ADD_11602

//ADD_6320 replaced by ADD_11602

//ADD_6330 replaced by ADD_11601

//ADD_6329 replaced by ADD_11602

//ADD_6328 replaced by ADD_11602

//ADD_6327 replaced by ADD_11602

//ADD_6326 replaced by ADD_11602

//ADD_6334 replaced by ADD_11602

//ADD_6333 replaced by ADD_11602

//ADD_6332 replaced by ADD_11602

//ADD_6331 replaced by ADD_11602

//BADD_1899 replaced by BADD_2824

//BADD_1898 replaced by BADD_2823

//BADD_1897 replaced by BADD_2822

//ADD_6336 replaced by ADD_11602

//ADD_6335 replaced by ADD_11602

//KaratsubaCore_659 replaced by KaratsubaCore_1437

//KaratsubaCore_658 replaced by KaratsubaCore_1438

//KaratsubaCore_657 replaced by KaratsubaCore_1437

//BADD_1903 replaced by BADD_2818

//BADD_1902 replaced by BADD_2820

//BADD_1901 replaced by BADD_2819

//BADD_1900 replaced by BADD_2818

//ADD_6338 replaced by ADD_8288

//ADD_6337 replaced by ADD_8288

//KaratsubaCore_662 replaced by KaratsubaCore_1438

//KaratsubaCore_661 replaced by KaratsubaCore_1435

//KaratsubaCore_660 replaced by KaratsubaCore_1438

//BADD_1906 replaced by BADD_2824

//BADD_1905 replaced by BADD_2823

//BADD_1904 replaced by BADD_2822

//ADD_6340 replaced by ADD_11602

//ADD_6339 replaced by ADD_11602

//KaratsubaCore_665 replaced by KaratsubaCore_1437

//KaratsubaCore_664 replaced by KaratsubaCore_1438

//KaratsubaCore_663 replaced by KaratsubaCore_1437

//ADD_6345 replaced by ADD_11595

//ADD_6344 replaced by ADD_11602

//ADD_6343 replaced by ADD_11602

//ADD_6342 replaced by ADD_11602

//ADD_6341 replaced by ADD_11602

//ADD_6350 replaced by ADD_11592

//ADD_6349 replaced by ADD_11602

//ADD_6348 replaced by ADD_11602

//ADD_6347 replaced by ADD_11602

//ADD_6346 replaced by ADD_11602

//ADD_6355 replaced by ADD_11592

//ADD_6354 replaced by ADD_11602

//ADD_6353 replaced by ADD_11602

//ADD_6352 replaced by ADD_11602

//ADD_6351 replaced by ADD_11602

//ADD_6360 replaced by ADD_11595

//ADD_6359 replaced by ADD_11602

//ADD_6358 replaced by ADD_11602

//ADD_6357 replaced by ADD_11602

//ADD_6356 replaced by ADD_11602

//BADD_1910 replaced by BADD_2818

//BADD_1909 replaced by BADD_2820

//BADD_1908 replaced by BADD_2819

//BADD_1907 replaced by BADD_2818

//ADD_6362 replaced by ADD_8288

//ADD_6361 replaced by ADD_8288

//KaratsubaCore_668 replaced by KaratsubaCore_1438

//KaratsubaCore_667 replaced by KaratsubaCore_1435

//KaratsubaCore_666 replaced by KaratsubaCore_1438

//BADD_1914 replaced by BADD_2807

//BADD_1913 replaced by BADD_2809

//BADD_1912 replaced by BADD_2808

//BADD_1911 replaced by BADD_2807

//ADD_6364 replaced by ADD_8267

//ADD_6363 replaced by ADD_8267

//KaratsubaCore_671 replaced by KaratsubaCore_1435

//KaratsubaCore_670 replaced by KaratsubaCore_1426

//KaratsubaCore_669 replaced by KaratsubaCore_1435

//BADD_1918 replaced by BADD_2818

//BADD_1917 replaced by BADD_2820

//BADD_1916 replaced by BADD_2819

//BADD_1915 replaced by BADD_2818

//ADD_6366 replaced by ADD_8288

//ADD_6365 replaced by ADD_8288

//KaratsubaCore_674 replaced by KaratsubaCore_1438

//KaratsubaCore_673 replaced by KaratsubaCore_1435

//KaratsubaCore_672 replaced by KaratsubaCore_1438

//ADD_6372 replaced by ADD_11602

//ADD_6371 replaced by ADD_11602

//ADD_6370 replaced by ADD_11602

//ADD_6369 replaced by ADD_11602

//ADD_6368 replaced by ADD_11602

//ADD_6367 replaced by ADD_11602

//ADD_6377 replaced by ADD_11601

//ADD_6376 replaced by ADD_11602

//ADD_6375 replaced by ADD_11602

//ADD_6374 replaced by ADD_11602

//ADD_6373 replaced by ADD_11602

//ADD_6381 replaced by ADD_11602

//ADD_6380 replaced by ADD_11602

//ADD_6379 replaced by ADD_11602

//ADD_6378 replaced by ADD_11602

//BADD_1921 replaced by BADD_2824

//BADD_1920 replaced by BADD_2823

//BADD_1919 replaced by BADD_2822

//ADD_6383 replaced by ADD_11602

//ADD_6382 replaced by ADD_11602

//KaratsubaCore_677 replaced by KaratsubaCore_1437

//KaratsubaCore_676 replaced by KaratsubaCore_1438

//KaratsubaCore_675 replaced by KaratsubaCore_1437

//BADD_1925 replaced by BADD_2818

//BADD_1924 replaced by BADD_2820

//BADD_1923 replaced by BADD_2819

//BADD_1922 replaced by BADD_2818

//ADD_6385 replaced by ADD_8288

//ADD_6384 replaced by ADD_8288

//KaratsubaCore_680 replaced by KaratsubaCore_1438

//KaratsubaCore_679 replaced by KaratsubaCore_1435

//KaratsubaCore_678 replaced by KaratsubaCore_1438

//BADD_1928 replaced by BADD_2824

//BADD_1927 replaced by BADD_2823

//BADD_1926 replaced by BADD_2822

//ADD_6387 replaced by ADD_11602

//ADD_6386 replaced by ADD_11602

//KaratsubaCore_683 replaced by KaratsubaCore_1437

//KaratsubaCore_682 replaced by KaratsubaCore_1438

//KaratsubaCore_681 replaced by KaratsubaCore_1437

//ADD_6393 replaced by ADD_11602

//ADD_6392 replaced by ADD_11602

//ADD_6391 replaced by ADD_11602

//ADD_6390 replaced by ADD_11602

//ADD_6389 replaced by ADD_11602

//ADD_6388 replaced by ADD_11602

//ADD_6398 replaced by ADD_11601

//ADD_6397 replaced by ADD_11602

//ADD_6396 replaced by ADD_11602

//ADD_6395 replaced by ADD_11602

//ADD_6394 replaced by ADD_11602

//ADD_6402 replaced by ADD_11602

//ADD_6401 replaced by ADD_11602

//ADD_6400 replaced by ADD_11602

//ADD_6399 replaced by ADD_11602

//BADD_1931 replaced by BADD_2824

//BADD_1930 replaced by BADD_2823

//BADD_1929 replaced by BADD_2822

//ADD_6404 replaced by ADD_11602

//ADD_6403 replaced by ADD_11602

//KaratsubaCore_686 replaced by KaratsubaCore_1437

//KaratsubaCore_685 replaced by KaratsubaCore_1438

//KaratsubaCore_684 replaced by KaratsubaCore_1437

//BADD_1935 replaced by BADD_2818

//BADD_1934 replaced by BADD_2820

//BADD_1933 replaced by BADD_2819

//BADD_1932 replaced by BADD_2818

//ADD_6406 replaced by ADD_8288

//ADD_6405 replaced by ADD_8288

//KaratsubaCore_689 replaced by KaratsubaCore_1438

//KaratsubaCore_688 replaced by KaratsubaCore_1435

//KaratsubaCore_687 replaced by KaratsubaCore_1438

//BADD_1938 replaced by BADD_2824

//BADD_1937 replaced by BADD_2823

//BADD_1936 replaced by BADD_2822

//ADD_6408 replaced by ADD_11602

//ADD_6407 replaced by ADD_11602

//KaratsubaCore_692 replaced by KaratsubaCore_1437

//KaratsubaCore_691 replaced by KaratsubaCore_1438

//KaratsubaCore_690 replaced by KaratsubaCore_1437

//ADD_6413 replaced by ADD_11595

//ADD_6412 replaced by ADD_11602

//ADD_6411 replaced by ADD_11602

//ADD_6410 replaced by ADD_11602

//ADD_6409 replaced by ADD_11602

//ADD_6418 replaced by ADD_11592

//ADD_6417 replaced by ADD_11602

//ADD_6416 replaced by ADD_11602

//ADD_6415 replaced by ADD_11602

//ADD_6414 replaced by ADD_11602

//ADD_6423 replaced by ADD_11592

//ADD_6422 replaced by ADD_11602

//ADD_6421 replaced by ADD_11602

//ADD_6420 replaced by ADD_11602

//ADD_6419 replaced by ADD_11602

//ADD_6428 replaced by ADD_11595

//ADD_6427 replaced by ADD_11602

//ADD_6426 replaced by ADD_11602

//ADD_6425 replaced by ADD_11602

//ADD_6424 replaced by ADD_11602

//BADD_1942 replaced by BADD_2818

//BADD_1941 replaced by BADD_2820

//BADD_1940 replaced by BADD_2819

//BADD_1939 replaced by BADD_2818

//ADD_6430 replaced by ADD_8288

//ADD_6429 replaced by ADD_8288

//KaratsubaCore_695 replaced by KaratsubaCore_1438

//KaratsubaCore_694 replaced by KaratsubaCore_1435

//KaratsubaCore_693 replaced by KaratsubaCore_1438

//BADD_1946 replaced by BADD_2807

//BADD_1945 replaced by BADD_2809

//BADD_1944 replaced by BADD_2808

//BADD_1943 replaced by BADD_2807

//ADD_6432 replaced by ADD_8267

//ADD_6431 replaced by ADD_8267

//KaratsubaCore_698 replaced by KaratsubaCore_1435

//KaratsubaCore_697 replaced by KaratsubaCore_1426

//KaratsubaCore_696 replaced by KaratsubaCore_1435

//BADD_1950 replaced by BADD_2818

//BADD_1949 replaced by BADD_2820

//BADD_1948 replaced by BADD_2819

//BADD_1947 replaced by BADD_2818

//ADD_6434 replaced by ADD_8288

//ADD_6433 replaced by ADD_8288

//KaratsubaCore_701 replaced by KaratsubaCore_1438

//KaratsubaCore_700 replaced by KaratsubaCore_1435

//KaratsubaCore_699 replaced by KaratsubaCore_1438

//ADD_6440 replaced by ADD_11602

//ADD_6439 replaced by ADD_11602

//ADD_6438 replaced by ADD_11602

//ADD_6437 replaced by ADD_11602

//ADD_6436 replaced by ADD_11602

//ADD_6435 replaced by ADD_11602

//ADD_6445 replaced by ADD_11601

//ADD_6444 replaced by ADD_11602

//ADD_6443 replaced by ADD_11602

//ADD_6442 replaced by ADD_11602

//ADD_6441 replaced by ADD_11602

//ADD_6449 replaced by ADD_11602

//ADD_6448 replaced by ADD_11602

//ADD_6447 replaced by ADD_11602

//ADD_6446 replaced by ADD_11602

//BADD_1953 replaced by BADD_2824

//BADD_1952 replaced by BADD_2823

//BADD_1951 replaced by BADD_2822

//ADD_6451 replaced by ADD_11602

//ADD_6450 replaced by ADD_11602

//KaratsubaCore_704 replaced by KaratsubaCore_1437

//KaratsubaCore_703 replaced by KaratsubaCore_1438

//KaratsubaCore_702 replaced by KaratsubaCore_1437

//BADD_1957 replaced by BADD_2818

//BADD_1956 replaced by BADD_2820

//BADD_1955 replaced by BADD_2819

//BADD_1954 replaced by BADD_2818

//ADD_6453 replaced by ADD_8288

//ADD_6452 replaced by ADD_8288

//KaratsubaCore_707 replaced by KaratsubaCore_1438

//KaratsubaCore_706 replaced by KaratsubaCore_1435

//KaratsubaCore_705 replaced by KaratsubaCore_1438

//BADD_1960 replaced by BADD_2824

//BADD_1959 replaced by BADD_2823

//BADD_1958 replaced by BADD_2822

//ADD_6455 replaced by ADD_11602

//ADD_6454 replaced by ADD_11602

//KaratsubaCore_710 replaced by KaratsubaCore_1437

//KaratsubaCore_709 replaced by KaratsubaCore_1438

//KaratsubaCore_708 replaced by KaratsubaCore_1437

//ADD_6461 replaced by ADD_11602

//ADD_6460 replaced by ADD_11602

//ADD_6459 replaced by ADD_11602

//ADD_6458 replaced by ADD_11602

//ADD_6457 replaced by ADD_11602

//ADD_6456 replaced by ADD_11602

//ADD_6466 replaced by ADD_11601

//ADD_6465 replaced by ADD_11602

//ADD_6464 replaced by ADD_11602

//ADD_6463 replaced by ADD_11602

//ADD_6462 replaced by ADD_11602

//ADD_6470 replaced by ADD_11602

//ADD_6469 replaced by ADD_11602

//ADD_6468 replaced by ADD_11602

//ADD_6467 replaced by ADD_11602

//BADD_1963 replaced by BADD_2824

//BADD_1962 replaced by BADD_2823

//BADD_1961 replaced by BADD_2822

//ADD_6472 replaced by ADD_11602

//ADD_6471 replaced by ADD_11602

//KaratsubaCore_713 replaced by KaratsubaCore_1437

//KaratsubaCore_712 replaced by KaratsubaCore_1438

//KaratsubaCore_711 replaced by KaratsubaCore_1437

//BADD_1967 replaced by BADD_2818

//BADD_1966 replaced by BADD_2820

//BADD_1965 replaced by BADD_2819

//BADD_1964 replaced by BADD_2818

//ADD_6474 replaced by ADD_8288

//ADD_6473 replaced by ADD_8288

//KaratsubaCore_716 replaced by KaratsubaCore_1438

//KaratsubaCore_715 replaced by KaratsubaCore_1435

//KaratsubaCore_714 replaced by KaratsubaCore_1438

//BADD_1970 replaced by BADD_2824

//BADD_1969 replaced by BADD_2823

//BADD_1968 replaced by BADD_2822

//ADD_6476 replaced by ADD_11602

//ADD_6475 replaced by ADD_11602

//KaratsubaCore_719 replaced by KaratsubaCore_1437

//KaratsubaCore_718 replaced by KaratsubaCore_1438

//KaratsubaCore_717 replaced by KaratsubaCore_1437

//ADD_6481 replaced by ADD_11595

//ADD_6480 replaced by ADD_11602

//ADD_6479 replaced by ADD_11602

//ADD_6478 replaced by ADD_11602

//ADD_6477 replaced by ADD_11602

//ADD_6486 replaced by ADD_11592

//ADD_6485 replaced by ADD_11602

//ADD_6484 replaced by ADD_11602

//ADD_6483 replaced by ADD_11602

//ADD_6482 replaced by ADD_11602

//ADD_6491 replaced by ADD_11592

//ADD_6490 replaced by ADD_11602

//ADD_6489 replaced by ADD_11602

//ADD_6488 replaced by ADD_11602

//ADD_6487 replaced by ADD_11602

//ADD_6496 replaced by ADD_11595

//ADD_6495 replaced by ADD_11602

//ADD_6494 replaced by ADD_11602

//ADD_6493 replaced by ADD_11602

//ADD_6492 replaced by ADD_11602

//BADD_1974 replaced by BADD_2818

//BADD_1973 replaced by BADD_2820

//BADD_1972 replaced by BADD_2819

//BADD_1971 replaced by BADD_2818

//ADD_6498 replaced by ADD_8288

//ADD_6497 replaced by ADD_8288

//KaratsubaCore_722 replaced by KaratsubaCore_1438

//KaratsubaCore_721 replaced by KaratsubaCore_1435

//KaratsubaCore_720 replaced by KaratsubaCore_1438

//BADD_1978 replaced by BADD_2807

//BADD_1977 replaced by BADD_2809

//BADD_1976 replaced by BADD_2808

//BADD_1975 replaced by BADD_2807

//ADD_6500 replaced by ADD_8267

//ADD_6499 replaced by ADD_8267

//KaratsubaCore_725 replaced by KaratsubaCore_1435

//KaratsubaCore_724 replaced by KaratsubaCore_1426

//KaratsubaCore_723 replaced by KaratsubaCore_1435

//BADD_1982 replaced by BADD_2818

//BADD_1981 replaced by BADD_2820

//BADD_1980 replaced by BADD_2819

//BADD_1979 replaced by BADD_2818

//ADD_6502 replaced by ADD_8288

//ADD_6501 replaced by ADD_8288

//KaratsubaCore_728 replaced by KaratsubaCore_1438

//KaratsubaCore_727 replaced by KaratsubaCore_1435

//KaratsubaCore_726 replaced by KaratsubaCore_1438

//ADD_6508 replaced by ADD_11602

//ADD_6507 replaced by ADD_11602

//ADD_6506 replaced by ADD_11602

//ADD_6505 replaced by ADD_11602

//ADD_6504 replaced by ADD_11602

//ADD_6503 replaced by ADD_11602

//ADD_6513 replaced by ADD_11601

//ADD_6512 replaced by ADD_11602

//ADD_6511 replaced by ADD_11602

//ADD_6510 replaced by ADD_11602

//ADD_6509 replaced by ADD_11602

//ADD_6517 replaced by ADD_11602

//ADD_6516 replaced by ADD_11602

//ADD_6515 replaced by ADD_11602

//ADD_6514 replaced by ADD_11602

//BADD_1985 replaced by BADD_2824

//BADD_1984 replaced by BADD_2823

//BADD_1983 replaced by BADD_2822

//ADD_6519 replaced by ADD_11602

//ADD_6518 replaced by ADD_11602

//KaratsubaCore_731 replaced by KaratsubaCore_1437

//KaratsubaCore_730 replaced by KaratsubaCore_1438

//KaratsubaCore_729 replaced by KaratsubaCore_1437

//BADD_1989 replaced by BADD_2818

//BADD_1988 replaced by BADD_2820

//BADD_1987 replaced by BADD_2819

//BADD_1986 replaced by BADD_2818

//ADD_6521 replaced by ADD_8288

//ADD_6520 replaced by ADD_8288

//KaratsubaCore_734 replaced by KaratsubaCore_1438

//KaratsubaCore_733 replaced by KaratsubaCore_1435

//KaratsubaCore_732 replaced by KaratsubaCore_1438

//BADD_1992 replaced by BADD_2824

//BADD_1991 replaced by BADD_2823

//BADD_1990 replaced by BADD_2822

//ADD_6523 replaced by ADD_11602

//ADD_6522 replaced by ADD_11602

//KaratsubaCore_737 replaced by KaratsubaCore_1437

//KaratsubaCore_736 replaced by KaratsubaCore_1438

//KaratsubaCore_735 replaced by KaratsubaCore_1437

//ADD_6529 replaced by ADD_11602

//ADD_6528 replaced by ADD_11602

//ADD_6527 replaced by ADD_11602

//ADD_6526 replaced by ADD_11602

//ADD_6525 replaced by ADD_11602

//ADD_6524 replaced by ADD_11602

//ADD_6534 replaced by ADD_11601

//ADD_6533 replaced by ADD_11602

//ADD_6532 replaced by ADD_11602

//ADD_6531 replaced by ADD_11602

//ADD_6530 replaced by ADD_11602

//ADD_6538 replaced by ADD_11602

//ADD_6537 replaced by ADD_11602

//ADD_6536 replaced by ADD_11602

//ADD_6535 replaced by ADD_11602

//BADD_1995 replaced by BADD_2824

//BADD_1994 replaced by BADD_2823

//BADD_1993 replaced by BADD_2822

//ADD_6540 replaced by ADD_11602

//ADD_6539 replaced by ADD_11602

//KaratsubaCore_740 replaced by KaratsubaCore_1437

//KaratsubaCore_739 replaced by KaratsubaCore_1438

//KaratsubaCore_738 replaced by KaratsubaCore_1437

//BADD_1999 replaced by BADD_2818

//BADD_1998 replaced by BADD_2820

//BADD_1997 replaced by BADD_2819

//BADD_1996 replaced by BADD_2818

//ADD_6542 replaced by ADD_8288

//ADD_6541 replaced by ADD_8288

//KaratsubaCore_743 replaced by KaratsubaCore_1438

//KaratsubaCore_742 replaced by KaratsubaCore_1435

//KaratsubaCore_741 replaced by KaratsubaCore_1438

//BADD_2002 replaced by BADD_2824

//BADD_2001 replaced by BADD_2823

//BADD_2000 replaced by BADD_2822

//ADD_6544 replaced by ADD_11602

//ADD_6543 replaced by ADD_11602

//KaratsubaCore_746 replaced by KaratsubaCore_1437

//KaratsubaCore_745 replaced by KaratsubaCore_1438

//KaratsubaCore_744 replaced by KaratsubaCore_1437

//ADD_6549 replaced by ADD_11595

//ADD_6548 replaced by ADD_11602

//ADD_6547 replaced by ADD_11602

//ADD_6546 replaced by ADD_11602

//ADD_6545 replaced by ADD_11602

//ADD_6554 replaced by ADD_11592

//ADD_6553 replaced by ADD_11602

//ADD_6552 replaced by ADD_11602

//ADD_6551 replaced by ADD_11602

//ADD_6550 replaced by ADD_11602

//ADD_6559 replaced by ADD_11592

//ADD_6558 replaced by ADD_11602

//ADD_6557 replaced by ADD_11602

//ADD_6556 replaced by ADD_11602

//ADD_6555 replaced by ADD_11602

//ADD_6564 replaced by ADD_11595

//ADD_6563 replaced by ADD_11602

//ADD_6562 replaced by ADD_11602

//ADD_6561 replaced by ADD_11602

//ADD_6560 replaced by ADD_11602

//BADD_2006 replaced by BADD_2818

//BADD_2005 replaced by BADD_2820

//BADD_2004 replaced by BADD_2819

//BADD_2003 replaced by BADD_2818

//ADD_6566 replaced by ADD_8288

//ADD_6565 replaced by ADD_8288

//KaratsubaCore_749 replaced by KaratsubaCore_1438

//KaratsubaCore_748 replaced by KaratsubaCore_1435

//KaratsubaCore_747 replaced by KaratsubaCore_1438

//BADD_2010 replaced by BADD_2807

//BADD_2009 replaced by BADD_2809

//BADD_2008 replaced by BADD_2808

//BADD_2007 replaced by BADD_2807

//ADD_6568 replaced by ADD_8267

//ADD_6567 replaced by ADD_8267

//KaratsubaCore_752 replaced by KaratsubaCore_1435

//KaratsubaCore_751 replaced by KaratsubaCore_1426

//KaratsubaCore_750 replaced by KaratsubaCore_1435

//BADD_2014 replaced by BADD_2818

//BADD_2013 replaced by BADD_2820

//BADD_2012 replaced by BADD_2819

//BADD_2011 replaced by BADD_2818

//ADD_6570 replaced by ADD_8288

//ADD_6569 replaced by ADD_8288

//KaratsubaCore_755 replaced by KaratsubaCore_1438

//KaratsubaCore_754 replaced by KaratsubaCore_1435

//KaratsubaCore_753 replaced by KaratsubaCore_1438

//ADD_6576 replaced by ADD_11602

//ADD_6575 replaced by ADD_11602

//ADD_6574 replaced by ADD_11602

//ADD_6573 replaced by ADD_11602

//ADD_6572 replaced by ADD_11602

//ADD_6571 replaced by ADD_11602

//ADD_6581 replaced by ADD_11601

//ADD_6580 replaced by ADD_11602

//ADD_6579 replaced by ADD_11602

//ADD_6578 replaced by ADD_11602

//ADD_6577 replaced by ADD_11602

//ADD_6585 replaced by ADD_11602

//ADD_6584 replaced by ADD_11602

//ADD_6583 replaced by ADD_11602

//ADD_6582 replaced by ADD_11602

//BADD_2017 replaced by BADD_2824

//BADD_2016 replaced by BADD_2823

//BADD_2015 replaced by BADD_2822

//ADD_6587 replaced by ADD_11602

//ADD_6586 replaced by ADD_11602

//KaratsubaCore_758 replaced by KaratsubaCore_1437

//KaratsubaCore_757 replaced by KaratsubaCore_1438

//KaratsubaCore_756 replaced by KaratsubaCore_1437

//BADD_2021 replaced by BADD_2818

//BADD_2020 replaced by BADD_2820

//BADD_2019 replaced by BADD_2819

//BADD_2018 replaced by BADD_2818

//ADD_6589 replaced by ADD_8288

//ADD_6588 replaced by ADD_8288

//KaratsubaCore_761 replaced by KaratsubaCore_1438

//KaratsubaCore_760 replaced by KaratsubaCore_1435

//KaratsubaCore_759 replaced by KaratsubaCore_1438

//BADD_2024 replaced by BADD_2824

//BADD_2023 replaced by BADD_2823

//BADD_2022 replaced by BADD_2822

//ADD_6591 replaced by ADD_11602

//ADD_6590 replaced by ADD_11602

//KaratsubaCore_764 replaced by KaratsubaCore_1437

//KaratsubaCore_763 replaced by KaratsubaCore_1438

//KaratsubaCore_762 replaced by KaratsubaCore_1437

//ADD_6597 replaced by ADD_11602

//ADD_6596 replaced by ADD_11602

//ADD_6595 replaced by ADD_11602

//ADD_6594 replaced by ADD_11602

//ADD_6593 replaced by ADD_11602

//ADD_6592 replaced by ADD_11602

//ADD_6602 replaced by ADD_11601

//ADD_6601 replaced by ADD_11602

//ADD_6600 replaced by ADD_11602

//ADD_6599 replaced by ADD_11602

//ADD_6598 replaced by ADD_11602

//ADD_6606 replaced by ADD_11602

//ADD_6605 replaced by ADD_11602

//ADD_6604 replaced by ADD_11602

//ADD_6603 replaced by ADD_11602

//BADD_2027 replaced by BADD_2824

//BADD_2026 replaced by BADD_2823

//BADD_2025 replaced by BADD_2822

//ADD_6608 replaced by ADD_11602

//ADD_6607 replaced by ADD_11602

//KaratsubaCore_767 replaced by KaratsubaCore_1437

//KaratsubaCore_766 replaced by KaratsubaCore_1438

//KaratsubaCore_765 replaced by KaratsubaCore_1437

//BADD_2031 replaced by BADD_2818

//BADD_2030 replaced by BADD_2820

//BADD_2029 replaced by BADD_2819

//BADD_2028 replaced by BADD_2818

//ADD_6610 replaced by ADD_8288

//ADD_6609 replaced by ADD_8288

//KaratsubaCore_770 replaced by KaratsubaCore_1438

//KaratsubaCore_769 replaced by KaratsubaCore_1435

//KaratsubaCore_768 replaced by KaratsubaCore_1438

//BADD_2034 replaced by BADD_2824

//BADD_2033 replaced by BADD_2823

//BADD_2032 replaced by BADD_2822

//ADD_6612 replaced by ADD_11602

//ADD_6611 replaced by ADD_11602

//KaratsubaCore_773 replaced by KaratsubaCore_1437

//KaratsubaCore_772 replaced by KaratsubaCore_1438

//KaratsubaCore_771 replaced by KaratsubaCore_1437

//ADD_6617 replaced by ADD_11595

//ADD_6616 replaced by ADD_11602

//ADD_6615 replaced by ADD_11602

//ADD_6614 replaced by ADD_11602

//ADD_6613 replaced by ADD_11602

//ADD_6622 replaced by ADD_11592

//ADD_6621 replaced by ADD_11602

//ADD_6620 replaced by ADD_11602

//ADD_6619 replaced by ADD_11602

//ADD_6618 replaced by ADD_11602

//ADD_6627 replaced by ADD_11592

//ADD_6626 replaced by ADD_11602

//ADD_6625 replaced by ADD_11602

//ADD_6624 replaced by ADD_11602

//ADD_6623 replaced by ADD_11602

//ADD_6632 replaced by ADD_11595

//ADD_6631 replaced by ADD_11602

//ADD_6630 replaced by ADD_11602

//ADD_6629 replaced by ADD_11602

//ADD_6628 replaced by ADD_11602

//BADD_2038 replaced by BADD_2818

//BADD_2037 replaced by BADD_2820

//BADD_2036 replaced by BADD_2819

//BADD_2035 replaced by BADD_2818

//ADD_6634 replaced by ADD_8288

//ADD_6633 replaced by ADD_8288

//KaratsubaCore_776 replaced by KaratsubaCore_1438

//KaratsubaCore_775 replaced by KaratsubaCore_1435

//KaratsubaCore_774 replaced by KaratsubaCore_1438

//BADD_2042 replaced by BADD_2807

//BADD_2041 replaced by BADD_2809

//BADD_2040 replaced by BADD_2808

//BADD_2039 replaced by BADD_2807

//ADD_6636 replaced by ADD_8267

//ADD_6635 replaced by ADD_8267

//KaratsubaCore_779 replaced by KaratsubaCore_1435

//KaratsubaCore_778 replaced by KaratsubaCore_1426

//KaratsubaCore_777 replaced by KaratsubaCore_1435

//BADD_2046 replaced by BADD_2818

//BADD_2045 replaced by BADD_2820

//BADD_2044 replaced by BADD_2819

//BADD_2043 replaced by BADD_2818

//ADD_6638 replaced by ADD_8288

//ADD_6637 replaced by ADD_8288

//KaratsubaCore_782 replaced by KaratsubaCore_1438

//KaratsubaCore_781 replaced by KaratsubaCore_1435

//KaratsubaCore_780 replaced by KaratsubaCore_1438

//ADD_6644 replaced by ADD_11602

//ADD_6643 replaced by ADD_11602

//ADD_6642 replaced by ADD_11602

//ADD_6641 replaced by ADD_11602

//ADD_6640 replaced by ADD_11602

//ADD_6639 replaced by ADD_11602

//ADD_6649 replaced by ADD_11601

//ADD_6648 replaced by ADD_11602

//ADD_6647 replaced by ADD_11602

//ADD_6646 replaced by ADD_11602

//ADD_6645 replaced by ADD_11602

//ADD_6653 replaced by ADD_11602

//ADD_6652 replaced by ADD_11602

//ADD_6651 replaced by ADD_11602

//ADD_6650 replaced by ADD_11602

//BADD_2049 replaced by BADD_2824

//BADD_2048 replaced by BADD_2823

//BADD_2047 replaced by BADD_2822

//ADD_6655 replaced by ADD_11602

//ADD_6654 replaced by ADD_11602

//KaratsubaCore_785 replaced by KaratsubaCore_1437

//KaratsubaCore_784 replaced by KaratsubaCore_1438

//KaratsubaCore_783 replaced by KaratsubaCore_1437

//BADD_2053 replaced by BADD_2818

//BADD_2052 replaced by BADD_2820

//BADD_2051 replaced by BADD_2819

//BADD_2050 replaced by BADD_2818

//ADD_6657 replaced by ADD_8288

//ADD_6656 replaced by ADD_8288

//KaratsubaCore_788 replaced by KaratsubaCore_1438

//KaratsubaCore_787 replaced by KaratsubaCore_1435

//KaratsubaCore_786 replaced by KaratsubaCore_1438

//BADD_2056 replaced by BADD_2824

//BADD_2055 replaced by BADD_2823

//BADD_2054 replaced by BADD_2822

//ADD_6659 replaced by ADD_11602

//ADD_6658 replaced by ADD_11602

//KaratsubaCore_791 replaced by KaratsubaCore_1437

//KaratsubaCore_790 replaced by KaratsubaCore_1438

//KaratsubaCore_789 replaced by KaratsubaCore_1437

//ADD_6665 replaced by ADD_11602

//ADD_6664 replaced by ADD_11602

//ADD_6663 replaced by ADD_11602

//ADD_6662 replaced by ADD_11602

//ADD_6661 replaced by ADD_11602

//ADD_6660 replaced by ADD_11602

//ADD_6670 replaced by ADD_11601

//ADD_6669 replaced by ADD_11602

//ADD_6668 replaced by ADD_11602

//ADD_6667 replaced by ADD_11602

//ADD_6666 replaced by ADD_11602

//ADD_6674 replaced by ADD_11602

//ADD_6673 replaced by ADD_11602

//ADD_6672 replaced by ADD_11602

//ADD_6671 replaced by ADD_11602

//BADD_2059 replaced by BADD_2824

//BADD_2058 replaced by BADD_2823

//BADD_2057 replaced by BADD_2822

//ADD_6676 replaced by ADD_11602

//ADD_6675 replaced by ADD_11602

//KaratsubaCore_794 replaced by KaratsubaCore_1437

//KaratsubaCore_793 replaced by KaratsubaCore_1438

//KaratsubaCore_792 replaced by KaratsubaCore_1437

//BADD_2063 replaced by BADD_2818

//BADD_2062 replaced by BADD_2820

//BADD_2061 replaced by BADD_2819

//BADD_2060 replaced by BADD_2818

//ADD_6678 replaced by ADD_8288

//ADD_6677 replaced by ADD_8288

//KaratsubaCore_797 replaced by KaratsubaCore_1438

//KaratsubaCore_796 replaced by KaratsubaCore_1435

//KaratsubaCore_795 replaced by KaratsubaCore_1438

//BADD_2066 replaced by BADD_2824

//BADD_2065 replaced by BADD_2823

//BADD_2064 replaced by BADD_2822

//ADD_6680 replaced by ADD_11602

//ADD_6679 replaced by ADD_11602

//KaratsubaCore_800 replaced by KaratsubaCore_1437

//KaratsubaCore_799 replaced by KaratsubaCore_1438

//KaratsubaCore_798 replaced by KaratsubaCore_1437

//ADD_6685 replaced by ADD_11595

//ADD_6684 replaced by ADD_11602

//ADD_6683 replaced by ADD_11602

//ADD_6682 replaced by ADD_11602

//ADD_6681 replaced by ADD_11602

//ADD_6690 replaced by ADD_11592

//ADD_6689 replaced by ADD_11602

//ADD_6688 replaced by ADD_11602

//ADD_6687 replaced by ADD_11602

//ADD_6686 replaced by ADD_11602

//ADD_6695 replaced by ADD_11592

//ADD_6694 replaced by ADD_11602

//ADD_6693 replaced by ADD_11602

//ADD_6692 replaced by ADD_11602

//ADD_6691 replaced by ADD_11602

//ADD_6700 replaced by ADD_11595

//ADD_6699 replaced by ADD_11602

//ADD_6698 replaced by ADD_11602

//ADD_6697 replaced by ADD_11602

//ADD_6696 replaced by ADD_11602

//BADD_2070 replaced by BADD_2818

//BADD_2069 replaced by BADD_2820

//BADD_2068 replaced by BADD_2819

//BADD_2067 replaced by BADD_2818

//ADD_6702 replaced by ADD_8288

//ADD_6701 replaced by ADD_8288

//KaratsubaCore_803 replaced by KaratsubaCore_1438

//KaratsubaCore_802 replaced by KaratsubaCore_1435

//KaratsubaCore_801 replaced by KaratsubaCore_1438

//BADD_2074 replaced by BADD_2807

//BADD_2073 replaced by BADD_2809

//BADD_2072 replaced by BADD_2808

//BADD_2071 replaced by BADD_2807

//ADD_6704 replaced by ADD_8267

//ADD_6703 replaced by ADD_8267

//KaratsubaCore_806 replaced by KaratsubaCore_1435

//KaratsubaCore_805 replaced by KaratsubaCore_1426

//KaratsubaCore_804 replaced by KaratsubaCore_1435

//BADD_2078 replaced by BADD_2818

//BADD_2077 replaced by BADD_2820

//BADD_2076 replaced by BADD_2819

//BADD_2075 replaced by BADD_2818

//ADD_6706 replaced by ADD_8288

//ADD_6705 replaced by ADD_8288

//KaratsubaCore_809 replaced by KaratsubaCore_1438

//KaratsubaCore_808 replaced by KaratsubaCore_1435

//KaratsubaCore_807 replaced by KaratsubaCore_1438

//ADD_6712 replaced by ADD_11602

//ADD_6711 replaced by ADD_11602

//ADD_6710 replaced by ADD_11602

//ADD_6709 replaced by ADD_11602

//ADD_6708 replaced by ADD_11602

//ADD_6707 replaced by ADD_11602

//ADD_6717 replaced by ADD_11601

//ADD_6716 replaced by ADD_11602

//ADD_6715 replaced by ADD_11602

//ADD_6714 replaced by ADD_11602

//ADD_6713 replaced by ADD_11602

//ADD_6721 replaced by ADD_11602

//ADD_6720 replaced by ADD_11602

//ADD_6719 replaced by ADD_11602

//ADD_6718 replaced by ADD_11602

//BADD_2081 replaced by BADD_2824

//BADD_2080 replaced by BADD_2823

//BADD_2079 replaced by BADD_2822

//ADD_6723 replaced by ADD_11602

//ADD_6722 replaced by ADD_11602

//KaratsubaCore_812 replaced by KaratsubaCore_1437

//KaratsubaCore_811 replaced by KaratsubaCore_1438

//KaratsubaCore_810 replaced by KaratsubaCore_1437

//BADD_2085 replaced by BADD_2818

//BADD_2084 replaced by BADD_2820

//BADD_2083 replaced by BADD_2819

//BADD_2082 replaced by BADD_2818

//ADD_6725 replaced by ADD_8288

//ADD_6724 replaced by ADD_8288

//KaratsubaCore_815 replaced by KaratsubaCore_1438

//KaratsubaCore_814 replaced by KaratsubaCore_1435

//KaratsubaCore_813 replaced by KaratsubaCore_1438

//BADD_2088 replaced by BADD_2824

//BADD_2087 replaced by BADD_2823

//BADD_2086 replaced by BADD_2822

//ADD_6727 replaced by ADD_11602

//ADD_6726 replaced by ADD_11602

//KaratsubaCore_818 replaced by KaratsubaCore_1437

//KaratsubaCore_817 replaced by KaratsubaCore_1438

//KaratsubaCore_816 replaced by KaratsubaCore_1437

//ADD_6733 replaced by ADD_11602

//ADD_6732 replaced by ADD_11602

//ADD_6731 replaced by ADD_11602

//ADD_6730 replaced by ADD_11602

//ADD_6729 replaced by ADD_11602

//ADD_6728 replaced by ADD_11602

//ADD_6738 replaced by ADD_11601

//ADD_6737 replaced by ADD_11602

//ADD_6736 replaced by ADD_11602

//ADD_6735 replaced by ADD_11602

//ADD_6734 replaced by ADD_11602

//ADD_6742 replaced by ADD_11602

//ADD_6741 replaced by ADD_11602

//ADD_6740 replaced by ADD_11602

//ADD_6739 replaced by ADD_11602

//BADD_2091 replaced by BADD_2824

//BADD_2090 replaced by BADD_2823

//BADD_2089 replaced by BADD_2822

//ADD_6744 replaced by ADD_11602

//ADD_6743 replaced by ADD_11602

//KaratsubaCore_821 replaced by KaratsubaCore_1437

//KaratsubaCore_820 replaced by KaratsubaCore_1438

//KaratsubaCore_819 replaced by KaratsubaCore_1437

//BADD_2095 replaced by BADD_2818

//BADD_2094 replaced by BADD_2820

//BADD_2093 replaced by BADD_2819

//BADD_2092 replaced by BADD_2818

//ADD_6746 replaced by ADD_8288

//ADD_6745 replaced by ADD_8288

//KaratsubaCore_824 replaced by KaratsubaCore_1438

//KaratsubaCore_823 replaced by KaratsubaCore_1435

//KaratsubaCore_822 replaced by KaratsubaCore_1438

//BADD_2098 replaced by BADD_2824

//BADD_2097 replaced by BADD_2823

//BADD_2096 replaced by BADD_2822

//ADD_6748 replaced by ADD_11602

//ADD_6747 replaced by ADD_11602

//KaratsubaCore_827 replaced by KaratsubaCore_1437

//KaratsubaCore_826 replaced by KaratsubaCore_1438

//KaratsubaCore_825 replaced by KaratsubaCore_1437

//ADD_6753 replaced by ADD_11595

//ADD_6752 replaced by ADD_11602

//ADD_6751 replaced by ADD_11602

//ADD_6750 replaced by ADD_11602

//ADD_6749 replaced by ADD_11602

//ADD_6758 replaced by ADD_11592

//ADD_6757 replaced by ADD_11602

//ADD_6756 replaced by ADD_11602

//ADD_6755 replaced by ADD_11602

//ADD_6754 replaced by ADD_11602

//ADD_6763 replaced by ADD_11592

//ADD_6762 replaced by ADD_11602

//ADD_6761 replaced by ADD_11602

//ADD_6760 replaced by ADD_11602

//ADD_6759 replaced by ADD_11602

//ADD_6768 replaced by ADD_11595

//ADD_6767 replaced by ADD_11602

//ADD_6766 replaced by ADD_11602

//ADD_6765 replaced by ADD_11602

//ADD_6764 replaced by ADD_11602

//BADD_2102 replaced by BADD_2818

//BADD_2101 replaced by BADD_2820

//BADD_2100 replaced by BADD_2819

//BADD_2099 replaced by BADD_2818

//ADD_6770 replaced by ADD_8288

//ADD_6769 replaced by ADD_8288

//KaratsubaCore_830 replaced by KaratsubaCore_1438

//KaratsubaCore_829 replaced by KaratsubaCore_1435

//KaratsubaCore_828 replaced by KaratsubaCore_1438

//BADD_2106 replaced by BADD_2807

//BADD_2105 replaced by BADD_2809

//BADD_2104 replaced by BADD_2808

//BADD_2103 replaced by BADD_2807

//ADD_6772 replaced by ADD_8267

//ADD_6771 replaced by ADD_8267

//KaratsubaCore_833 replaced by KaratsubaCore_1435

//KaratsubaCore_832 replaced by KaratsubaCore_1426

//KaratsubaCore_831 replaced by KaratsubaCore_1435

//BADD_2110 replaced by BADD_2818

//BADD_2109 replaced by BADD_2820

//BADD_2108 replaced by BADD_2819

//BADD_2107 replaced by BADD_2818

//ADD_6774 replaced by ADD_8288

//ADD_6773 replaced by ADD_8288

//KaratsubaCore_836 replaced by KaratsubaCore_1438

//KaratsubaCore_835 replaced by KaratsubaCore_1435

//KaratsubaCore_834 replaced by KaratsubaCore_1438

//ADD_6780 replaced by ADD_11602

//ADD_6779 replaced by ADD_11602

//ADD_6778 replaced by ADD_11602

//ADD_6777 replaced by ADD_11602

//ADD_6776 replaced by ADD_11602

//ADD_6775 replaced by ADD_11602

//ADD_6785 replaced by ADD_11601

//ADD_6784 replaced by ADD_11602

//ADD_6783 replaced by ADD_11602

//ADD_6782 replaced by ADD_11602

//ADD_6781 replaced by ADD_11602

//ADD_6789 replaced by ADD_11602

//ADD_6788 replaced by ADD_11602

//ADD_6787 replaced by ADD_11602

//ADD_6786 replaced by ADD_11602

//BADD_2113 replaced by BADD_2824

//BADD_2112 replaced by BADD_2823

//BADD_2111 replaced by BADD_2822

//ADD_6791 replaced by ADD_11602

//ADD_6790 replaced by ADD_11602

//KaratsubaCore_839 replaced by KaratsubaCore_1437

//KaratsubaCore_838 replaced by KaratsubaCore_1438

//KaratsubaCore_837 replaced by KaratsubaCore_1437

//BADD_2117 replaced by BADD_2818

//BADD_2116 replaced by BADD_2820

//BADD_2115 replaced by BADD_2819

//BADD_2114 replaced by BADD_2818

//ADD_6793 replaced by ADD_8288

//ADD_6792 replaced by ADD_8288

//KaratsubaCore_842 replaced by KaratsubaCore_1438

//KaratsubaCore_841 replaced by KaratsubaCore_1435

//KaratsubaCore_840 replaced by KaratsubaCore_1438

//BADD_2120 replaced by BADD_2824

//BADD_2119 replaced by BADD_2823

//BADD_2118 replaced by BADD_2822

//ADD_6795 replaced by ADD_11602

//ADD_6794 replaced by ADD_11602

//KaratsubaCore_845 replaced by KaratsubaCore_1437

//KaratsubaCore_844 replaced by KaratsubaCore_1438

//KaratsubaCore_843 replaced by KaratsubaCore_1437

//ADD_6801 replaced by ADD_11602

//ADD_6800 replaced by ADD_11602

//ADD_6799 replaced by ADD_11602

//ADD_6798 replaced by ADD_11602

//ADD_6797 replaced by ADD_11602

//ADD_6796 replaced by ADD_11602

//ADD_6806 replaced by ADD_11601

//ADD_6805 replaced by ADD_11602

//ADD_6804 replaced by ADD_11602

//ADD_6803 replaced by ADD_11602

//ADD_6802 replaced by ADD_11602

//ADD_6810 replaced by ADD_11602

//ADD_6809 replaced by ADD_11602

//ADD_6808 replaced by ADD_11602

//ADD_6807 replaced by ADD_11602

//BADD_2123 replaced by BADD_2824

//BADD_2122 replaced by BADD_2823

//BADD_2121 replaced by BADD_2822

//ADD_6812 replaced by ADD_11602

//ADD_6811 replaced by ADD_11602

//KaratsubaCore_848 replaced by KaratsubaCore_1437

//KaratsubaCore_847 replaced by KaratsubaCore_1438

//KaratsubaCore_846 replaced by KaratsubaCore_1437

//BADD_2127 replaced by BADD_2818

//BADD_2126 replaced by BADD_2820

//BADD_2125 replaced by BADD_2819

//BADD_2124 replaced by BADD_2818

//ADD_6814 replaced by ADD_8288

//ADD_6813 replaced by ADD_8288

//KaratsubaCore_851 replaced by KaratsubaCore_1438

//KaratsubaCore_850 replaced by KaratsubaCore_1435

//KaratsubaCore_849 replaced by KaratsubaCore_1438

//BADD_2130 replaced by BADD_2824

//BADD_2129 replaced by BADD_2823

//BADD_2128 replaced by BADD_2822

//ADD_6816 replaced by ADD_11602

//ADD_6815 replaced by ADD_11602

//KaratsubaCore_854 replaced by KaratsubaCore_1437

//KaratsubaCore_853 replaced by KaratsubaCore_1438

//KaratsubaCore_852 replaced by KaratsubaCore_1437

//ADD_6821 replaced by ADD_11595

//ADD_6820 replaced by ADD_11602

//ADD_6819 replaced by ADD_11602

//ADD_6818 replaced by ADD_11602

//ADD_6817 replaced by ADD_11602

//ADD_6826 replaced by ADD_11592

//ADD_6825 replaced by ADD_11602

//ADD_6824 replaced by ADD_11602

//ADD_6823 replaced by ADD_11602

//ADD_6822 replaced by ADD_11602

//ADD_6831 replaced by ADD_11592

//ADD_6830 replaced by ADD_11602

//ADD_6829 replaced by ADD_11602

//ADD_6828 replaced by ADD_11602

//ADD_6827 replaced by ADD_11602

//ADD_6836 replaced by ADD_11595

//ADD_6835 replaced by ADD_11602

//ADD_6834 replaced by ADD_11602

//ADD_6833 replaced by ADD_11602

//ADD_6832 replaced by ADD_11602

//BADD_2134 replaced by BADD_2818

//BADD_2133 replaced by BADD_2820

//BADD_2132 replaced by BADD_2819

//BADD_2131 replaced by BADD_2818

//ADD_6838 replaced by ADD_8288

//ADD_6837 replaced by ADD_8288

//KaratsubaCore_857 replaced by KaratsubaCore_1438

//KaratsubaCore_856 replaced by KaratsubaCore_1435

//KaratsubaCore_855 replaced by KaratsubaCore_1438

//BADD_2138 replaced by BADD_2807

//BADD_2137 replaced by BADD_2809

//BADD_2136 replaced by BADD_2808

//BADD_2135 replaced by BADD_2807

//ADD_6840 replaced by ADD_8267

//ADD_6839 replaced by ADD_8267

//KaratsubaCore_860 replaced by KaratsubaCore_1435

//KaratsubaCore_859 replaced by KaratsubaCore_1426

//KaratsubaCore_858 replaced by KaratsubaCore_1435

//BADD_2142 replaced by BADD_2818

//BADD_2141 replaced by BADD_2820

//BADD_2140 replaced by BADD_2819

//BADD_2139 replaced by BADD_2818

//ADD_6842 replaced by ADD_8288

//ADD_6841 replaced by ADD_8288

//KaratsubaCore_863 replaced by KaratsubaCore_1438

//KaratsubaCore_862 replaced by KaratsubaCore_1435

//KaratsubaCore_861 replaced by KaratsubaCore_1438

//ADD_6848 replaced by ADD_11602

//ADD_6847 replaced by ADD_11602

//ADD_6846 replaced by ADD_11602

//ADD_6845 replaced by ADD_11602

//ADD_6844 replaced by ADD_11602

//ADD_6843 replaced by ADD_11602

//ADD_6853 replaced by ADD_11601

//ADD_6852 replaced by ADD_11602

//ADD_6851 replaced by ADD_11602

//ADD_6850 replaced by ADD_11602

//ADD_6849 replaced by ADD_11602

//ADD_6857 replaced by ADD_11602

//ADD_6856 replaced by ADD_11602

//ADD_6855 replaced by ADD_11602

//ADD_6854 replaced by ADD_11602

//BADD_2145 replaced by BADD_2824

//BADD_2144 replaced by BADD_2823

//BADD_2143 replaced by BADD_2822

//ADD_6859 replaced by ADD_11602

//ADD_6858 replaced by ADD_11602

//KaratsubaCore_866 replaced by KaratsubaCore_1437

//KaratsubaCore_865 replaced by KaratsubaCore_1438

//KaratsubaCore_864 replaced by KaratsubaCore_1437

//BADD_2149 replaced by BADD_2818

//BADD_2148 replaced by BADD_2820

//BADD_2147 replaced by BADD_2819

//BADD_2146 replaced by BADD_2818

//ADD_6861 replaced by ADD_8288

//ADD_6860 replaced by ADD_8288

//KaratsubaCore_869 replaced by KaratsubaCore_1438

//KaratsubaCore_868 replaced by KaratsubaCore_1435

//KaratsubaCore_867 replaced by KaratsubaCore_1438

//BADD_2152 replaced by BADD_2824

//BADD_2151 replaced by BADD_2823

//BADD_2150 replaced by BADD_2822

//ADD_6863 replaced by ADD_11602

//ADD_6862 replaced by ADD_11602

//KaratsubaCore_872 replaced by KaratsubaCore_1437

//KaratsubaCore_871 replaced by KaratsubaCore_1438

//KaratsubaCore_870 replaced by KaratsubaCore_1437

//ADD_6869 replaced by ADD_11602

//ADD_6868 replaced by ADD_11602

//ADD_6867 replaced by ADD_11602

//ADD_6866 replaced by ADD_11602

//ADD_6865 replaced by ADD_11602

//ADD_6864 replaced by ADD_11602

//ADD_6874 replaced by ADD_11601

//ADD_6873 replaced by ADD_11602

//ADD_6872 replaced by ADD_11602

//ADD_6871 replaced by ADD_11602

//ADD_6870 replaced by ADD_11602

//ADD_6878 replaced by ADD_11602

//ADD_6877 replaced by ADD_11602

//ADD_6876 replaced by ADD_11602

//ADD_6875 replaced by ADD_11602

//BADD_2155 replaced by BADD_2824

//BADD_2154 replaced by BADD_2823

//BADD_2153 replaced by BADD_2822

//ADD_6880 replaced by ADD_11602

//ADD_6879 replaced by ADD_11602

//KaratsubaCore_875 replaced by KaratsubaCore_1437

//KaratsubaCore_874 replaced by KaratsubaCore_1438

//KaratsubaCore_873 replaced by KaratsubaCore_1437

//BADD_2159 replaced by BADD_2818

//BADD_2158 replaced by BADD_2820

//BADD_2157 replaced by BADD_2819

//BADD_2156 replaced by BADD_2818

//ADD_6882 replaced by ADD_8288

//ADD_6881 replaced by ADD_8288

//KaratsubaCore_878 replaced by KaratsubaCore_1438

//KaratsubaCore_877 replaced by KaratsubaCore_1435

//KaratsubaCore_876 replaced by KaratsubaCore_1438

//BADD_2162 replaced by BADD_2824

//BADD_2161 replaced by BADD_2823

//BADD_2160 replaced by BADD_2822

//ADD_6884 replaced by ADD_11602

//ADD_6883 replaced by ADD_11602

//KaratsubaCore_881 replaced by KaratsubaCore_1437

//KaratsubaCore_880 replaced by KaratsubaCore_1438

//KaratsubaCore_879 replaced by KaratsubaCore_1437

//ADD_6889 replaced by ADD_11595

//ADD_6888 replaced by ADD_11602

//ADD_6887 replaced by ADD_11602

//ADD_6886 replaced by ADD_11602

//ADD_6885 replaced by ADD_11602

//ADD_6894 replaced by ADD_11592

//ADD_6893 replaced by ADD_11602

//ADD_6892 replaced by ADD_11602

//ADD_6891 replaced by ADD_11602

//ADD_6890 replaced by ADD_11602

//ADD_6899 replaced by ADD_11592

//ADD_6898 replaced by ADD_11602

//ADD_6897 replaced by ADD_11602

//ADD_6896 replaced by ADD_11602

//ADD_6895 replaced by ADD_11602

//ADD_6904 replaced by ADD_11595

//ADD_6903 replaced by ADD_11602

//ADD_6902 replaced by ADD_11602

//ADD_6901 replaced by ADD_11602

//ADD_6900 replaced by ADD_11602

//BADD_2166 replaced by BADD_2818

//BADD_2165 replaced by BADD_2820

//BADD_2164 replaced by BADD_2819

//BADD_2163 replaced by BADD_2818

//ADD_6906 replaced by ADD_8288

//ADD_6905 replaced by ADD_8288

//KaratsubaCore_884 replaced by KaratsubaCore_1438

//KaratsubaCore_883 replaced by KaratsubaCore_1435

//KaratsubaCore_882 replaced by KaratsubaCore_1438

//BADD_2170 replaced by BADD_2807

//BADD_2169 replaced by BADD_2809

//BADD_2168 replaced by BADD_2808

//BADD_2167 replaced by BADD_2807

//ADD_6908 replaced by ADD_8267

//ADD_6907 replaced by ADD_8267

//KaratsubaCore_887 replaced by KaratsubaCore_1435

//KaratsubaCore_886 replaced by KaratsubaCore_1426

//KaratsubaCore_885 replaced by KaratsubaCore_1435

//BADD_2174 replaced by BADD_2818

//BADD_2173 replaced by BADD_2820

//BADD_2172 replaced by BADD_2819

//BADD_2171 replaced by BADD_2818

//ADD_6910 replaced by ADD_8288

//ADD_6909 replaced by ADD_8288

//KaratsubaCore_890 replaced by KaratsubaCore_1438

//KaratsubaCore_889 replaced by KaratsubaCore_1435

//KaratsubaCore_888 replaced by KaratsubaCore_1438

//ADD_6916 replaced by ADD_11602

//ADD_6915 replaced by ADD_11602

//ADD_6914 replaced by ADD_11602

//ADD_6913 replaced by ADD_11602

//ADD_6912 replaced by ADD_11602

//ADD_6911 replaced by ADD_11602

//ADD_6921 replaced by ADD_11601

//ADD_6920 replaced by ADD_11602

//ADD_6919 replaced by ADD_11602

//ADD_6918 replaced by ADD_11602

//ADD_6917 replaced by ADD_11602

//ADD_6925 replaced by ADD_11602

//ADD_6924 replaced by ADD_11602

//ADD_6923 replaced by ADD_11602

//ADD_6922 replaced by ADD_11602

//BADD_2177 replaced by BADD_2824

//BADD_2176 replaced by BADD_2823

//BADD_2175 replaced by BADD_2822

//ADD_6927 replaced by ADD_11602

//ADD_6926 replaced by ADD_11602

//KaratsubaCore_893 replaced by KaratsubaCore_1437

//KaratsubaCore_892 replaced by KaratsubaCore_1438

//KaratsubaCore_891 replaced by KaratsubaCore_1437

//BADD_2181 replaced by BADD_2818

//BADD_2180 replaced by BADD_2820

//BADD_2179 replaced by BADD_2819

//BADD_2178 replaced by BADD_2818

//ADD_6929 replaced by ADD_8288

//ADD_6928 replaced by ADD_8288

//KaratsubaCore_896 replaced by KaratsubaCore_1438

//KaratsubaCore_895 replaced by KaratsubaCore_1435

//KaratsubaCore_894 replaced by KaratsubaCore_1438

//BADD_2184 replaced by BADD_2824

//BADD_2183 replaced by BADD_2823

//BADD_2182 replaced by BADD_2822

//ADD_6931 replaced by ADD_11602

//ADD_6930 replaced by ADD_11602

//KaratsubaCore_899 replaced by KaratsubaCore_1437

//KaratsubaCore_898 replaced by KaratsubaCore_1438

//KaratsubaCore_897 replaced by KaratsubaCore_1437

//ADD_6937 replaced by ADD_11602

//ADD_6936 replaced by ADD_11602

//ADD_6935 replaced by ADD_11602

//ADD_6934 replaced by ADD_11602

//ADD_6933 replaced by ADD_11602

//ADD_6932 replaced by ADD_11602

//ADD_6942 replaced by ADD_11601

//ADD_6941 replaced by ADD_11602

//ADD_6940 replaced by ADD_11602

//ADD_6939 replaced by ADD_11602

//ADD_6938 replaced by ADD_11602

//ADD_6946 replaced by ADD_11602

//ADD_6945 replaced by ADD_11602

//ADD_6944 replaced by ADD_11602

//ADD_6943 replaced by ADD_11602

//BADD_2187 replaced by BADD_2824

//BADD_2186 replaced by BADD_2823

//BADD_2185 replaced by BADD_2822

//ADD_6948 replaced by ADD_11602

//ADD_6947 replaced by ADD_11602

//KaratsubaCore_902 replaced by KaratsubaCore_1437

//KaratsubaCore_901 replaced by KaratsubaCore_1438

//KaratsubaCore_900 replaced by KaratsubaCore_1437

//BADD_2191 replaced by BADD_2818

//BADD_2190 replaced by BADD_2820

//BADD_2189 replaced by BADD_2819

//BADD_2188 replaced by BADD_2818

//ADD_6950 replaced by ADD_8288

//ADD_6949 replaced by ADD_8288

//KaratsubaCore_905 replaced by KaratsubaCore_1438

//KaratsubaCore_904 replaced by KaratsubaCore_1435

//KaratsubaCore_903 replaced by KaratsubaCore_1438

//BADD_2194 replaced by BADD_2824

//BADD_2193 replaced by BADD_2823

//BADD_2192 replaced by BADD_2822

//ADD_6952 replaced by ADD_11602

//ADD_6951 replaced by ADD_11602

//KaratsubaCore_908 replaced by KaratsubaCore_1437

//KaratsubaCore_907 replaced by KaratsubaCore_1438

//KaratsubaCore_906 replaced by KaratsubaCore_1437

//ADD_6957 replaced by ADD_11595

//ADD_6956 replaced by ADD_11602

//ADD_6955 replaced by ADD_11602

//ADD_6954 replaced by ADD_11602

//ADD_6953 replaced by ADD_11602

//ADD_6962 replaced by ADD_11592

//ADD_6961 replaced by ADD_11602

//ADD_6960 replaced by ADD_11602

//ADD_6959 replaced by ADD_11602

//ADD_6958 replaced by ADD_11602

//ADD_6967 replaced by ADD_11592

//ADD_6966 replaced by ADD_11602

//ADD_6965 replaced by ADD_11602

//ADD_6964 replaced by ADD_11602

//ADD_6963 replaced by ADD_11602

//ADD_6972 replaced by ADD_11595

//ADD_6971 replaced by ADD_11602

//ADD_6970 replaced by ADD_11602

//ADD_6969 replaced by ADD_11602

//ADD_6968 replaced by ADD_11602

//BADD_2198 replaced by BADD_2818

//BADD_2197 replaced by BADD_2820

//BADD_2196 replaced by BADD_2819

//BADD_2195 replaced by BADD_2818

//ADD_6974 replaced by ADD_8288

//ADD_6973 replaced by ADD_8288

//KaratsubaCore_911 replaced by KaratsubaCore_1438

//KaratsubaCore_910 replaced by KaratsubaCore_1435

//KaratsubaCore_909 replaced by KaratsubaCore_1438

//BADD_2202 replaced by BADD_2807

//BADD_2201 replaced by BADD_2809

//BADD_2200 replaced by BADD_2808

//BADD_2199 replaced by BADD_2807

//ADD_6976 replaced by ADD_8267

//ADD_6975 replaced by ADD_8267

//KaratsubaCore_914 replaced by KaratsubaCore_1435

//KaratsubaCore_913 replaced by KaratsubaCore_1426

//KaratsubaCore_912 replaced by KaratsubaCore_1435

//BADD_2206 replaced by BADD_2818

//BADD_2205 replaced by BADD_2820

//BADD_2204 replaced by BADD_2819

//BADD_2203 replaced by BADD_2818

//ADD_6978 replaced by ADD_8288

//ADD_6977 replaced by ADD_8288

//KaratsubaCore_917 replaced by KaratsubaCore_1438

//KaratsubaCore_916 replaced by KaratsubaCore_1435

//KaratsubaCore_915 replaced by KaratsubaCore_1438

//ADD_6984 replaced by ADD_11602

//ADD_6983 replaced by ADD_11602

//ADD_6982 replaced by ADD_11602

//ADD_6981 replaced by ADD_11602

//ADD_6980 replaced by ADD_11602

//ADD_6979 replaced by ADD_11602

//ADD_6989 replaced by ADD_11601

//ADD_6988 replaced by ADD_11602

//ADD_6987 replaced by ADD_11602

//ADD_6986 replaced by ADD_11602

//ADD_6985 replaced by ADD_11602

//ADD_6993 replaced by ADD_11602

//ADD_6992 replaced by ADD_11602

//ADD_6991 replaced by ADD_11602

//ADD_6990 replaced by ADD_11602

//BADD_2209 replaced by BADD_2824

//BADD_2208 replaced by BADD_2823

//BADD_2207 replaced by BADD_2822

//ADD_6995 replaced by ADD_11602

//ADD_6994 replaced by ADD_11602

//KaratsubaCore_920 replaced by KaratsubaCore_1437

//KaratsubaCore_919 replaced by KaratsubaCore_1438

//KaratsubaCore_918 replaced by KaratsubaCore_1437

//BADD_2213 replaced by BADD_2818

//BADD_2212 replaced by BADD_2820

//BADD_2211 replaced by BADD_2819

//BADD_2210 replaced by BADD_2818

//ADD_6997 replaced by ADD_8288

//ADD_6996 replaced by ADD_8288

//KaratsubaCore_923 replaced by KaratsubaCore_1438

//KaratsubaCore_922 replaced by KaratsubaCore_1435

//KaratsubaCore_921 replaced by KaratsubaCore_1438

//BADD_2216 replaced by BADD_2824

//BADD_2215 replaced by BADD_2823

//BADD_2214 replaced by BADD_2822

//ADD_6999 replaced by ADD_11602

//ADD_6998 replaced by ADD_11602

//KaratsubaCore_926 replaced by KaratsubaCore_1437

//KaratsubaCore_925 replaced by KaratsubaCore_1438

//KaratsubaCore_924 replaced by KaratsubaCore_1437

//ADD_7005 replaced by ADD_11602

//ADD_7004 replaced by ADD_11602

//ADD_7003 replaced by ADD_11602

//ADD_7002 replaced by ADD_11602

//ADD_7001 replaced by ADD_11602

//ADD_7000 replaced by ADD_11602

//ADD_7010 replaced by ADD_11601

//ADD_7009 replaced by ADD_11602

//ADD_7008 replaced by ADD_11602

//ADD_7007 replaced by ADD_11602

//ADD_7006 replaced by ADD_11602

//ADD_7014 replaced by ADD_11602

//ADD_7013 replaced by ADD_11602

//ADD_7012 replaced by ADD_11602

//ADD_7011 replaced by ADD_11602

//BADD_2219 replaced by BADD_2824

//BADD_2218 replaced by BADD_2823

//BADD_2217 replaced by BADD_2822

//ADD_7016 replaced by ADD_11602

//ADD_7015 replaced by ADD_11602

//KaratsubaCore_929 replaced by KaratsubaCore_1437

//KaratsubaCore_928 replaced by KaratsubaCore_1438

//KaratsubaCore_927 replaced by KaratsubaCore_1437

//BADD_2223 replaced by BADD_2818

//BADD_2222 replaced by BADD_2820

//BADD_2221 replaced by BADD_2819

//BADD_2220 replaced by BADD_2818

//ADD_7018 replaced by ADD_8288

//ADD_7017 replaced by ADD_8288

//KaratsubaCore_932 replaced by KaratsubaCore_1438

//KaratsubaCore_931 replaced by KaratsubaCore_1435

//KaratsubaCore_930 replaced by KaratsubaCore_1438

//BADD_2226 replaced by BADD_2824

//BADD_2225 replaced by BADD_2823

//BADD_2224 replaced by BADD_2822

//ADD_7020 replaced by ADD_11602

//ADD_7019 replaced by ADD_11602

//KaratsubaCore_935 replaced by KaratsubaCore_1437

//KaratsubaCore_934 replaced by KaratsubaCore_1438

//KaratsubaCore_933 replaced by KaratsubaCore_1437

//ADD_7025 replaced by ADD_11595

//ADD_7024 replaced by ADD_11602

//ADD_7023 replaced by ADD_11602

//ADD_7022 replaced by ADD_11602

//ADD_7021 replaced by ADD_11602

//ADD_7030 replaced by ADD_11592

//ADD_7029 replaced by ADD_11602

//ADD_7028 replaced by ADD_11602

//ADD_7027 replaced by ADD_11602

//ADD_7026 replaced by ADD_11602

//ADD_7035 replaced by ADD_11592

//ADD_7034 replaced by ADD_11602

//ADD_7033 replaced by ADD_11602

//ADD_7032 replaced by ADD_11602

//ADD_7031 replaced by ADD_11602

//ADD_7040 replaced by ADD_11595

//ADD_7039 replaced by ADD_11602

//ADD_7038 replaced by ADD_11602

//ADD_7037 replaced by ADD_11602

//ADD_7036 replaced by ADD_11602

//BADD_2230 replaced by BADD_2818

//BADD_2229 replaced by BADD_2820

//BADD_2228 replaced by BADD_2819

//BADD_2227 replaced by BADD_2818

//ADD_7042 replaced by ADD_8288

//ADD_7041 replaced by ADD_8288

//KaratsubaCore_938 replaced by KaratsubaCore_1438

//KaratsubaCore_937 replaced by KaratsubaCore_1435

//KaratsubaCore_936 replaced by KaratsubaCore_1438

//BADD_2234 replaced by BADD_2807

//BADD_2233 replaced by BADD_2809

//BADD_2232 replaced by BADD_2808

//BADD_2231 replaced by BADD_2807

//ADD_7044 replaced by ADD_8267

//ADD_7043 replaced by ADD_8267

//KaratsubaCore_941 replaced by KaratsubaCore_1435

//KaratsubaCore_940 replaced by KaratsubaCore_1426

//KaratsubaCore_939 replaced by KaratsubaCore_1435

//BADD_2238 replaced by BADD_2818

//BADD_2237 replaced by BADD_2820

//BADD_2236 replaced by BADD_2819

//BADD_2235 replaced by BADD_2818

//ADD_7046 replaced by ADD_8288

//ADD_7045 replaced by ADD_8288

//KaratsubaCore_944 replaced by KaratsubaCore_1438

//KaratsubaCore_943 replaced by KaratsubaCore_1435

//KaratsubaCore_942 replaced by KaratsubaCore_1438

//ADD_7052 replaced by ADD_11602

//ADD_7051 replaced by ADD_11602

//ADD_7050 replaced by ADD_11602

//ADD_7049 replaced by ADD_11602

//ADD_7048 replaced by ADD_11602

//ADD_7047 replaced by ADD_11602

//ADD_7057 replaced by ADD_11601

//ADD_7056 replaced by ADD_11602

//ADD_7055 replaced by ADD_11602

//ADD_7054 replaced by ADD_11602

//ADD_7053 replaced by ADD_11602

//ADD_7061 replaced by ADD_11602

//ADD_7060 replaced by ADD_11602

//ADD_7059 replaced by ADD_11602

//ADD_7058 replaced by ADD_11602

//BADD_2241 replaced by BADD_2824

//BADD_2240 replaced by BADD_2823

//BADD_2239 replaced by BADD_2822

//ADD_7063 replaced by ADD_11602

//ADD_7062 replaced by ADD_11602

//KaratsubaCore_947 replaced by KaratsubaCore_1437

//KaratsubaCore_946 replaced by KaratsubaCore_1438

//KaratsubaCore_945 replaced by KaratsubaCore_1437

//BADD_2245 replaced by BADD_2818

//BADD_2244 replaced by BADD_2820

//BADD_2243 replaced by BADD_2819

//BADD_2242 replaced by BADD_2818

//ADD_7065 replaced by ADD_8288

//ADD_7064 replaced by ADD_8288

//KaratsubaCore_950 replaced by KaratsubaCore_1438

//KaratsubaCore_949 replaced by KaratsubaCore_1435

//KaratsubaCore_948 replaced by KaratsubaCore_1438

//BADD_2248 replaced by BADD_2824

//BADD_2247 replaced by BADD_2823

//BADD_2246 replaced by BADD_2822

//ADD_7067 replaced by ADD_11602

//ADD_7066 replaced by ADD_11602

//KaratsubaCore_953 replaced by KaratsubaCore_1437

//KaratsubaCore_952 replaced by KaratsubaCore_1438

//KaratsubaCore_951 replaced by KaratsubaCore_1437

//ADD_7073 replaced by ADD_11602

//ADD_7072 replaced by ADD_11602

//ADD_7071 replaced by ADD_11602

//ADD_7070 replaced by ADD_11602

//ADD_7069 replaced by ADD_11602

//ADD_7068 replaced by ADD_11602

//ADD_7078 replaced by ADD_11601

//ADD_7077 replaced by ADD_11602

//ADD_7076 replaced by ADD_11602

//ADD_7075 replaced by ADD_11602

//ADD_7074 replaced by ADD_11602

//ADD_7082 replaced by ADD_11602

//ADD_7081 replaced by ADD_11602

//ADD_7080 replaced by ADD_11602

//ADD_7079 replaced by ADD_11602

//BADD_2251 replaced by BADD_2824

//BADD_2250 replaced by BADD_2823

//BADD_2249 replaced by BADD_2822

//ADD_7084 replaced by ADD_11602

//ADD_7083 replaced by ADD_11602

//KaratsubaCore_956 replaced by KaratsubaCore_1437

//KaratsubaCore_955 replaced by KaratsubaCore_1438

//KaratsubaCore_954 replaced by KaratsubaCore_1437

//BADD_2255 replaced by BADD_2818

//BADD_2254 replaced by BADD_2820

//BADD_2253 replaced by BADD_2819

//BADD_2252 replaced by BADD_2818

//ADD_7086 replaced by ADD_8288

//ADD_7085 replaced by ADD_8288

//KaratsubaCore_959 replaced by KaratsubaCore_1438

//KaratsubaCore_958 replaced by KaratsubaCore_1435

//KaratsubaCore_957 replaced by KaratsubaCore_1438

//BADD_2258 replaced by BADD_2824

//BADD_2257 replaced by BADD_2823

//BADD_2256 replaced by BADD_2822

//ADD_7088 replaced by ADD_11602

//ADD_7087 replaced by ADD_11602

//KaratsubaCore_962 replaced by KaratsubaCore_1437

//KaratsubaCore_961 replaced by KaratsubaCore_1438

//KaratsubaCore_960 replaced by KaratsubaCore_1437

//ADD_7093 replaced by ADD_11595

//ADD_7092 replaced by ADD_11602

//ADD_7091 replaced by ADD_11602

//ADD_7090 replaced by ADD_11602

//ADD_7089 replaced by ADD_11602

//ADD_7098 replaced by ADD_11592

//ADD_7097 replaced by ADD_11602

//ADD_7096 replaced by ADD_11602

//ADD_7095 replaced by ADD_11602

//ADD_7094 replaced by ADD_11602

//ADD_7103 replaced by ADD_11592

//ADD_7102 replaced by ADD_11602

//ADD_7101 replaced by ADD_11602

//ADD_7100 replaced by ADD_11602

//ADD_7099 replaced by ADD_11602

//ADD_7108 replaced by ADD_11595

//ADD_7107 replaced by ADD_11602

//ADD_7106 replaced by ADD_11602

//ADD_7105 replaced by ADD_11602

//ADD_7104 replaced by ADD_11602

//BADD_2262 replaced by BADD_2818

//BADD_2261 replaced by BADD_2820

//BADD_2260 replaced by BADD_2819

//BADD_2259 replaced by BADD_2818

//ADD_7110 replaced by ADD_8288

//ADD_7109 replaced by ADD_8288

//KaratsubaCore_965 replaced by KaratsubaCore_1438

//KaratsubaCore_964 replaced by KaratsubaCore_1435

//KaratsubaCore_963 replaced by KaratsubaCore_1438

//BADD_2266 replaced by BADD_2807

//BADD_2265 replaced by BADD_2809

//BADD_2264 replaced by BADD_2808

//BADD_2263 replaced by BADD_2807

//ADD_7112 replaced by ADD_8267

//ADD_7111 replaced by ADD_8267

//KaratsubaCore_968 replaced by KaratsubaCore_1435

//KaratsubaCore_967 replaced by KaratsubaCore_1426

//KaratsubaCore_966 replaced by KaratsubaCore_1435

//BADD_2270 replaced by BADD_2818

//BADD_2269 replaced by BADD_2820

//BADD_2268 replaced by BADD_2819

//BADD_2267 replaced by BADD_2818

//ADD_7114 replaced by ADD_8288

//ADD_7113 replaced by ADD_8288

//KaratsubaCore_971 replaced by KaratsubaCore_1438

//KaratsubaCore_970 replaced by KaratsubaCore_1435

//KaratsubaCore_969 replaced by KaratsubaCore_1438

//ADD_7120 replaced by ADD_11602

//ADD_7119 replaced by ADD_11602

//ADD_7118 replaced by ADD_11602

//ADD_7117 replaced by ADD_11602

//ADD_7116 replaced by ADD_11602

//ADD_7115 replaced by ADD_11602

//ADD_7125 replaced by ADD_11601

//ADD_7124 replaced by ADD_11602

//ADD_7123 replaced by ADD_11602

//ADD_7122 replaced by ADD_11602

//ADD_7121 replaced by ADD_11602

//ADD_7129 replaced by ADD_11602

//ADD_7128 replaced by ADD_11602

//ADD_7127 replaced by ADD_11602

//ADD_7126 replaced by ADD_11602

//BADD_2273 replaced by BADD_2824

//BADD_2272 replaced by BADD_2823

//BADD_2271 replaced by BADD_2822

//ADD_7131 replaced by ADD_11602

//ADD_7130 replaced by ADD_11602

//KaratsubaCore_974 replaced by KaratsubaCore_1437

//KaratsubaCore_973 replaced by KaratsubaCore_1438

//KaratsubaCore_972 replaced by KaratsubaCore_1437

//BADD_2277 replaced by BADD_2818

//BADD_2276 replaced by BADD_2820

//BADD_2275 replaced by BADD_2819

//BADD_2274 replaced by BADD_2818

//ADD_7133 replaced by ADD_8288

//ADD_7132 replaced by ADD_8288

//KaratsubaCore_977 replaced by KaratsubaCore_1438

//KaratsubaCore_976 replaced by KaratsubaCore_1435

//KaratsubaCore_975 replaced by KaratsubaCore_1438

//BADD_2280 replaced by BADD_2824

//BADD_2279 replaced by BADD_2823

//BADD_2278 replaced by BADD_2822

//ADD_7135 replaced by ADD_11602

//ADD_7134 replaced by ADD_11602

//KaratsubaCore_980 replaced by KaratsubaCore_1437

//KaratsubaCore_979 replaced by KaratsubaCore_1438

//KaratsubaCore_978 replaced by KaratsubaCore_1437

//ADD_7141 replaced by ADD_11602

//ADD_7140 replaced by ADD_11602

//ADD_7139 replaced by ADD_11602

//ADD_7138 replaced by ADD_11602

//ADD_7137 replaced by ADD_11602

//ADD_7136 replaced by ADD_11602

//ADD_7146 replaced by ADD_11601

//ADD_7145 replaced by ADD_11602

//ADD_7144 replaced by ADD_11602

//ADD_7143 replaced by ADD_11602

//ADD_7142 replaced by ADD_11602

//ADD_7150 replaced by ADD_11602

//ADD_7149 replaced by ADD_11602

//ADD_7148 replaced by ADD_11602

//ADD_7147 replaced by ADD_11602

//BADD_2283 replaced by BADD_2824

//BADD_2282 replaced by BADD_2823

//BADD_2281 replaced by BADD_2822

//ADD_7152 replaced by ADD_11602

//ADD_7151 replaced by ADD_11602

//KaratsubaCore_983 replaced by KaratsubaCore_1437

//KaratsubaCore_982 replaced by KaratsubaCore_1438

//KaratsubaCore_981 replaced by KaratsubaCore_1437

//BADD_2287 replaced by BADD_2818

//BADD_2286 replaced by BADD_2820

//BADD_2285 replaced by BADD_2819

//BADD_2284 replaced by BADD_2818

//ADD_7154 replaced by ADD_8288

//ADD_7153 replaced by ADD_8288

//KaratsubaCore_986 replaced by KaratsubaCore_1438

//KaratsubaCore_985 replaced by KaratsubaCore_1435

//KaratsubaCore_984 replaced by KaratsubaCore_1438

//BADD_2290 replaced by BADD_2824

//BADD_2289 replaced by BADD_2823

//BADD_2288 replaced by BADD_2822

//ADD_7156 replaced by ADD_11602

//ADD_7155 replaced by ADD_11602

//KaratsubaCore_989 replaced by KaratsubaCore_1437

//KaratsubaCore_988 replaced by KaratsubaCore_1438

//KaratsubaCore_987 replaced by KaratsubaCore_1437

//ADD_7161 replaced by ADD_11595

//ADD_7160 replaced by ADD_11602

//ADD_7159 replaced by ADD_11602

//ADD_7158 replaced by ADD_11602

//ADD_7157 replaced by ADD_11602

//ADD_7166 replaced by ADD_11592

//ADD_7165 replaced by ADD_11602

//ADD_7164 replaced by ADD_11602

//ADD_7163 replaced by ADD_11602

//ADD_7162 replaced by ADD_11602

//ADD_7171 replaced by ADD_11592

//ADD_7170 replaced by ADD_11602

//ADD_7169 replaced by ADD_11602

//ADD_7168 replaced by ADD_11602

//ADD_7167 replaced by ADD_11602

//ADD_7176 replaced by ADD_11595

//ADD_7175 replaced by ADD_11602

//ADD_7174 replaced by ADD_11602

//ADD_7173 replaced by ADD_11602

//ADD_7172 replaced by ADD_11602

//BADD_2294 replaced by BADD_2818

//BADD_2293 replaced by BADD_2820

//BADD_2292 replaced by BADD_2819

//BADD_2291 replaced by BADD_2818

//ADD_7178 replaced by ADD_8288

//ADD_7177 replaced by ADD_8288

//KaratsubaCore_992 replaced by KaratsubaCore_1438

//KaratsubaCore_991 replaced by KaratsubaCore_1435

//KaratsubaCore_990 replaced by KaratsubaCore_1438

//BADD_2298 replaced by BADD_2807

//BADD_2297 replaced by BADD_2809

//BADD_2296 replaced by BADD_2808

//BADD_2295 replaced by BADD_2807

//ADD_7180 replaced by ADD_8267

//ADD_7179 replaced by ADD_8267

//KaratsubaCore_995 replaced by KaratsubaCore_1435

//KaratsubaCore_994 replaced by KaratsubaCore_1426

//KaratsubaCore_993 replaced by KaratsubaCore_1435

//BADD_2302 replaced by BADD_2818

//BADD_2301 replaced by BADD_2820

//BADD_2300 replaced by BADD_2819

//BADD_2299 replaced by BADD_2818

//ADD_7182 replaced by ADD_8288

//ADD_7181 replaced by ADD_8288

//KaratsubaCore_998 replaced by KaratsubaCore_1438

//KaratsubaCore_997 replaced by KaratsubaCore_1435

//KaratsubaCore_996 replaced by KaratsubaCore_1438

//ADD_7188 replaced by ADD_11602

//ADD_7187 replaced by ADD_11602

//ADD_7186 replaced by ADD_11602

//ADD_7185 replaced by ADD_11602

//ADD_7184 replaced by ADD_11602

//ADD_7183 replaced by ADD_11602

//ADD_7193 replaced by ADD_11601

//ADD_7192 replaced by ADD_11602

//ADD_7191 replaced by ADD_11602

//ADD_7190 replaced by ADD_11602

//ADD_7189 replaced by ADD_11602

//ADD_7197 replaced by ADD_11602

//ADD_7196 replaced by ADD_11602

//ADD_7195 replaced by ADD_11602

//ADD_7194 replaced by ADD_11602

//BADD_2305 replaced by BADD_2824

//BADD_2304 replaced by BADD_2823

//BADD_2303 replaced by BADD_2822

//ADD_7199 replaced by ADD_11602

//ADD_7198 replaced by ADD_11602

//KaratsubaCore_1001 replaced by KaratsubaCore_1437

//KaratsubaCore_1000 replaced by KaratsubaCore_1438

//KaratsubaCore_999 replaced by KaratsubaCore_1437

//BADD_2309 replaced by BADD_2818

//BADD_2308 replaced by BADD_2820

//BADD_2307 replaced by BADD_2819

//BADD_2306 replaced by BADD_2818

//ADD_7201 replaced by ADD_8288

//ADD_7200 replaced by ADD_8288

//KaratsubaCore_1004 replaced by KaratsubaCore_1438

//KaratsubaCore_1003 replaced by KaratsubaCore_1435

//KaratsubaCore_1002 replaced by KaratsubaCore_1438

//BADD_2312 replaced by BADD_2824

//BADD_2311 replaced by BADD_2823

//BADD_2310 replaced by BADD_2822

//ADD_7203 replaced by ADD_11602

//ADD_7202 replaced by ADD_11602

//KaratsubaCore_1007 replaced by KaratsubaCore_1437

//KaratsubaCore_1006 replaced by KaratsubaCore_1438

//KaratsubaCore_1005 replaced by KaratsubaCore_1437

//ADD_7209 replaced by ADD_11602

//ADD_7208 replaced by ADD_11602

//ADD_7207 replaced by ADD_11602

//ADD_7206 replaced by ADD_11602

//ADD_7205 replaced by ADD_11602

//ADD_7204 replaced by ADD_11602

//ADD_7214 replaced by ADD_11601

//ADD_7213 replaced by ADD_11602

//ADD_7212 replaced by ADD_11602

//ADD_7211 replaced by ADD_11602

//ADD_7210 replaced by ADD_11602

//ADD_7218 replaced by ADD_11602

//ADD_7217 replaced by ADD_11602

//ADD_7216 replaced by ADD_11602

//ADD_7215 replaced by ADD_11602

//BADD_2315 replaced by BADD_2824

//BADD_2314 replaced by BADD_2823

//BADD_2313 replaced by BADD_2822

//ADD_7220 replaced by ADD_11602

//ADD_7219 replaced by ADD_11602

//KaratsubaCore_1010 replaced by KaratsubaCore_1437

//KaratsubaCore_1009 replaced by KaratsubaCore_1438

//KaratsubaCore_1008 replaced by KaratsubaCore_1437

//BADD_2319 replaced by BADD_2818

//BADD_2318 replaced by BADD_2820

//BADD_2317 replaced by BADD_2819

//BADD_2316 replaced by BADD_2818

//ADD_7222 replaced by ADD_8288

//ADD_7221 replaced by ADD_8288

//KaratsubaCore_1013 replaced by KaratsubaCore_1438

//KaratsubaCore_1012 replaced by KaratsubaCore_1435

//KaratsubaCore_1011 replaced by KaratsubaCore_1438

//BADD_2322 replaced by BADD_2824

//BADD_2321 replaced by BADD_2823

//BADD_2320 replaced by BADD_2822

//ADD_7224 replaced by ADD_11602

//ADD_7223 replaced by ADD_11602

//KaratsubaCore_1016 replaced by KaratsubaCore_1437

//KaratsubaCore_1015 replaced by KaratsubaCore_1438

//KaratsubaCore_1014 replaced by KaratsubaCore_1437

//ADD_7229 replaced by ADD_11595

//ADD_7228 replaced by ADD_11602

//ADD_7227 replaced by ADD_11602

//ADD_7226 replaced by ADD_11602

//ADD_7225 replaced by ADD_11602

//ADD_7234 replaced by ADD_11592

//ADD_7233 replaced by ADD_11602

//ADD_7232 replaced by ADD_11602

//ADD_7231 replaced by ADD_11602

//ADD_7230 replaced by ADD_11602

//ADD_7239 replaced by ADD_11592

//ADD_7238 replaced by ADD_11602

//ADD_7237 replaced by ADD_11602

//ADD_7236 replaced by ADD_11602

//ADD_7235 replaced by ADD_11602

//ADD_7244 replaced by ADD_11595

//ADD_7243 replaced by ADD_11602

//ADD_7242 replaced by ADD_11602

//ADD_7241 replaced by ADD_11602

//ADD_7240 replaced by ADD_11602

//BADD_2326 replaced by BADD_2818

//BADD_2325 replaced by BADD_2820

//BADD_2324 replaced by BADD_2819

//BADD_2323 replaced by BADD_2818

//ADD_7246 replaced by ADD_8288

//ADD_7245 replaced by ADD_8288

//KaratsubaCore_1019 replaced by KaratsubaCore_1438

//KaratsubaCore_1018 replaced by KaratsubaCore_1435

//KaratsubaCore_1017 replaced by KaratsubaCore_1438

//BADD_2330 replaced by BADD_2807

//BADD_2329 replaced by BADD_2809

//BADD_2328 replaced by BADD_2808

//BADD_2327 replaced by BADD_2807

//ADD_7248 replaced by ADD_8267

//ADD_7247 replaced by ADD_8267

//KaratsubaCore_1022 replaced by KaratsubaCore_1435

//KaratsubaCore_1021 replaced by KaratsubaCore_1426

//KaratsubaCore_1020 replaced by KaratsubaCore_1435

//BADD_2334 replaced by BADD_2818

//BADD_2333 replaced by BADD_2820

//BADD_2332 replaced by BADD_2819

//BADD_2331 replaced by BADD_2818

//ADD_7250 replaced by ADD_8288

//ADD_7249 replaced by ADD_8288

//KaratsubaCore_1025 replaced by KaratsubaCore_1438

//KaratsubaCore_1024 replaced by KaratsubaCore_1435

//KaratsubaCore_1023 replaced by KaratsubaCore_1438

//ADD_7256 replaced by ADD_11602

//ADD_7255 replaced by ADD_11602

//ADD_7254 replaced by ADD_11602

//ADD_7253 replaced by ADD_11602

//ADD_7252 replaced by ADD_11602

//ADD_7251 replaced by ADD_11602

//ADD_7261 replaced by ADD_11601

//ADD_7260 replaced by ADD_11602

//ADD_7259 replaced by ADD_11602

//ADD_7258 replaced by ADD_11602

//ADD_7257 replaced by ADD_11602

//ADD_7265 replaced by ADD_11602

//ADD_7264 replaced by ADD_11602

//ADD_7263 replaced by ADD_11602

//ADD_7262 replaced by ADD_11602

//BADD_2337 replaced by BADD_2824

//BADD_2336 replaced by BADD_2823

//BADD_2335 replaced by BADD_2822

//ADD_7267 replaced by ADD_11602

//ADD_7266 replaced by ADD_11602

//KaratsubaCore_1028 replaced by KaratsubaCore_1437

//KaratsubaCore_1027 replaced by KaratsubaCore_1438

//KaratsubaCore_1026 replaced by KaratsubaCore_1437

//BADD_2341 replaced by BADD_2818

//BADD_2340 replaced by BADD_2820

//BADD_2339 replaced by BADD_2819

//BADD_2338 replaced by BADD_2818

//ADD_7269 replaced by ADD_8288

//ADD_7268 replaced by ADD_8288

//KaratsubaCore_1031 replaced by KaratsubaCore_1438

//KaratsubaCore_1030 replaced by KaratsubaCore_1435

//KaratsubaCore_1029 replaced by KaratsubaCore_1438

//BADD_2344 replaced by BADD_2824

//BADD_2343 replaced by BADD_2823

//BADD_2342 replaced by BADD_2822

//ADD_7271 replaced by ADD_11602

//ADD_7270 replaced by ADD_11602

//KaratsubaCore_1034 replaced by KaratsubaCore_1437

//KaratsubaCore_1033 replaced by KaratsubaCore_1438

//KaratsubaCore_1032 replaced by KaratsubaCore_1437

//ADD_7277 replaced by ADD_11602

//ADD_7276 replaced by ADD_11602

//ADD_7275 replaced by ADD_11602

//ADD_7274 replaced by ADD_11602

//ADD_7273 replaced by ADD_11602

//ADD_7272 replaced by ADD_11602

//ADD_7282 replaced by ADD_11601

//ADD_7281 replaced by ADD_11602

//ADD_7280 replaced by ADD_11602

//ADD_7279 replaced by ADD_11602

//ADD_7278 replaced by ADD_11602

//ADD_7286 replaced by ADD_11602

//ADD_7285 replaced by ADD_11602

//ADD_7284 replaced by ADD_11602

//ADD_7283 replaced by ADD_11602

//BADD_2347 replaced by BADD_2824

//BADD_2346 replaced by BADD_2823

//BADD_2345 replaced by BADD_2822

//ADD_7288 replaced by ADD_11602

//ADD_7287 replaced by ADD_11602

//KaratsubaCore_1037 replaced by KaratsubaCore_1437

//KaratsubaCore_1036 replaced by KaratsubaCore_1438

//KaratsubaCore_1035 replaced by KaratsubaCore_1437

//BADD_2351 replaced by BADD_2818

//BADD_2350 replaced by BADD_2820

//BADD_2349 replaced by BADD_2819

//BADD_2348 replaced by BADD_2818

//ADD_7290 replaced by ADD_8288

//ADD_7289 replaced by ADD_8288

//KaratsubaCore_1040 replaced by KaratsubaCore_1438

//KaratsubaCore_1039 replaced by KaratsubaCore_1435

//KaratsubaCore_1038 replaced by KaratsubaCore_1438

//BADD_2354 replaced by BADD_2824

//BADD_2353 replaced by BADD_2823

//BADD_2352 replaced by BADD_2822

//ADD_7292 replaced by ADD_11602

//ADD_7291 replaced by ADD_11602

//KaratsubaCore_1043 replaced by KaratsubaCore_1437

//KaratsubaCore_1042 replaced by KaratsubaCore_1438

//KaratsubaCore_1041 replaced by KaratsubaCore_1437

//ADD_7297 replaced by ADD_11595

//ADD_7296 replaced by ADD_11602

//ADD_7295 replaced by ADD_11602

//ADD_7294 replaced by ADD_11602

//ADD_7293 replaced by ADD_11602

//ADD_7302 replaced by ADD_11592

//ADD_7301 replaced by ADD_11602

//ADD_7300 replaced by ADD_11602

//ADD_7299 replaced by ADD_11602

//ADD_7298 replaced by ADD_11602

//ADD_7307 replaced by ADD_11592

//ADD_7306 replaced by ADD_11602

//ADD_7305 replaced by ADD_11602

//ADD_7304 replaced by ADD_11602

//ADD_7303 replaced by ADD_11602

//ADD_7312 replaced by ADD_11595

//ADD_7311 replaced by ADD_11602

//ADD_7310 replaced by ADD_11602

//ADD_7309 replaced by ADD_11602

//ADD_7308 replaced by ADD_11602

//BADD_2358 replaced by BADD_2818

//BADD_2357 replaced by BADD_2820

//BADD_2356 replaced by BADD_2819

//BADD_2355 replaced by BADD_2818

//ADD_7314 replaced by ADD_8288

//ADD_7313 replaced by ADD_8288

//KaratsubaCore_1046 replaced by KaratsubaCore_1438

//KaratsubaCore_1045 replaced by KaratsubaCore_1435

//KaratsubaCore_1044 replaced by KaratsubaCore_1438

//BADD_2362 replaced by BADD_2807

//BADD_2361 replaced by BADD_2809

//BADD_2360 replaced by BADD_2808

//BADD_2359 replaced by BADD_2807

//ADD_7316 replaced by ADD_8267

//ADD_7315 replaced by ADD_8267

//KaratsubaCore_1049 replaced by KaratsubaCore_1435

//KaratsubaCore_1048 replaced by KaratsubaCore_1426

//KaratsubaCore_1047 replaced by KaratsubaCore_1435

//BADD_2366 replaced by BADD_2818

//BADD_2365 replaced by BADD_2820

//BADD_2364 replaced by BADD_2819

//BADD_2363 replaced by BADD_2818

//ADD_7318 replaced by ADD_8288

//ADD_7317 replaced by ADD_8288

//KaratsubaCore_1052 replaced by KaratsubaCore_1438

//KaratsubaCore_1051 replaced by KaratsubaCore_1435

//KaratsubaCore_1050 replaced by KaratsubaCore_1438

//ADD_7324 replaced by ADD_11602

//ADD_7323 replaced by ADD_11602

//ADD_7322 replaced by ADD_11602

//ADD_7321 replaced by ADD_11602

//ADD_7320 replaced by ADD_11602

//ADD_7319 replaced by ADD_11602

//ADD_7329 replaced by ADD_11601

//ADD_7328 replaced by ADD_11602

//ADD_7327 replaced by ADD_11602

//ADD_7326 replaced by ADD_11602

//ADD_7325 replaced by ADD_11602

//ADD_7333 replaced by ADD_11602

//ADD_7332 replaced by ADD_11602

//ADD_7331 replaced by ADD_11602

//ADD_7330 replaced by ADD_11602

//BADD_2369 replaced by BADD_2824

//BADD_2368 replaced by BADD_2823

//BADD_2367 replaced by BADD_2822

//ADD_7335 replaced by ADD_11602

//ADD_7334 replaced by ADD_11602

//KaratsubaCore_1055 replaced by KaratsubaCore_1437

//KaratsubaCore_1054 replaced by KaratsubaCore_1438

//KaratsubaCore_1053 replaced by KaratsubaCore_1437

//BADD_2373 replaced by BADD_2818

//BADD_2372 replaced by BADD_2820

//BADD_2371 replaced by BADD_2819

//BADD_2370 replaced by BADD_2818

//ADD_7337 replaced by ADD_8288

//ADD_7336 replaced by ADD_8288

//KaratsubaCore_1058 replaced by KaratsubaCore_1438

//KaratsubaCore_1057 replaced by KaratsubaCore_1435

//KaratsubaCore_1056 replaced by KaratsubaCore_1438

//BADD_2376 replaced by BADD_2824

//BADD_2375 replaced by BADD_2823

//BADD_2374 replaced by BADD_2822

//ADD_7339 replaced by ADD_11602

//ADD_7338 replaced by ADD_11602

//KaratsubaCore_1061 replaced by KaratsubaCore_1437

//KaratsubaCore_1060 replaced by KaratsubaCore_1438

//KaratsubaCore_1059 replaced by KaratsubaCore_1437

//ADD_7345 replaced by ADD_11602

//ADD_7344 replaced by ADD_11602

//ADD_7343 replaced by ADD_11602

//ADD_7342 replaced by ADD_11602

//ADD_7341 replaced by ADD_11602

//ADD_7340 replaced by ADD_11602

//ADD_7350 replaced by ADD_11601

//ADD_7349 replaced by ADD_11602

//ADD_7348 replaced by ADD_11602

//ADD_7347 replaced by ADD_11602

//ADD_7346 replaced by ADD_11602

//ADD_7354 replaced by ADD_11602

//ADD_7353 replaced by ADD_11602

//ADD_7352 replaced by ADD_11602

//ADD_7351 replaced by ADD_11602

//BADD_2379 replaced by BADD_2824

//BADD_2378 replaced by BADD_2823

//BADD_2377 replaced by BADD_2822

//ADD_7356 replaced by ADD_11602

//ADD_7355 replaced by ADD_11602

//KaratsubaCore_1064 replaced by KaratsubaCore_1437

//KaratsubaCore_1063 replaced by KaratsubaCore_1438

//KaratsubaCore_1062 replaced by KaratsubaCore_1437

//BADD_2383 replaced by BADD_2818

//BADD_2382 replaced by BADD_2820

//BADD_2381 replaced by BADD_2819

//BADD_2380 replaced by BADD_2818

//ADD_7358 replaced by ADD_8288

//ADD_7357 replaced by ADD_8288

//KaratsubaCore_1067 replaced by KaratsubaCore_1438

//KaratsubaCore_1066 replaced by KaratsubaCore_1435

//KaratsubaCore_1065 replaced by KaratsubaCore_1438

//BADD_2386 replaced by BADD_2824

//BADD_2385 replaced by BADD_2823

//BADD_2384 replaced by BADD_2822

//ADD_7360 replaced by ADD_11602

//ADD_7359 replaced by ADD_11602

//KaratsubaCore_1070 replaced by KaratsubaCore_1437

//KaratsubaCore_1069 replaced by KaratsubaCore_1438

//KaratsubaCore_1068 replaced by KaratsubaCore_1437

//ADD_7365 replaced by ADD_11595

//ADD_7364 replaced by ADD_11602

//ADD_7363 replaced by ADD_11602

//ADD_7362 replaced by ADD_11602

//ADD_7361 replaced by ADD_11602

//ADD_7370 replaced by ADD_11592

//ADD_7369 replaced by ADD_11602

//ADD_7368 replaced by ADD_11602

//ADD_7367 replaced by ADD_11602

//ADD_7366 replaced by ADD_11602

//ADD_7375 replaced by ADD_11592

//ADD_7374 replaced by ADD_11602

//ADD_7373 replaced by ADD_11602

//ADD_7372 replaced by ADD_11602

//ADD_7371 replaced by ADD_11602

//ADD_7380 replaced by ADD_11595

//ADD_7379 replaced by ADD_11602

//ADD_7378 replaced by ADD_11602

//ADD_7377 replaced by ADD_11602

//ADD_7376 replaced by ADD_11602

//BADD_2390 replaced by BADD_2818

//BADD_2389 replaced by BADD_2820

//BADD_2388 replaced by BADD_2819

//BADD_2387 replaced by BADD_2818

//ADD_7382 replaced by ADD_8288

//ADD_7381 replaced by ADD_8288

//KaratsubaCore_1073 replaced by KaratsubaCore_1438

//KaratsubaCore_1072 replaced by KaratsubaCore_1435

//KaratsubaCore_1071 replaced by KaratsubaCore_1438

//BADD_2394 replaced by BADD_2807

//BADD_2393 replaced by BADD_2809

//BADD_2392 replaced by BADD_2808

//BADD_2391 replaced by BADD_2807

//ADD_7384 replaced by ADD_8267

//ADD_7383 replaced by ADD_8267

//KaratsubaCore_1076 replaced by KaratsubaCore_1435

//KaratsubaCore_1075 replaced by KaratsubaCore_1426

//KaratsubaCore_1074 replaced by KaratsubaCore_1435

//BADD_2398 replaced by BADD_2818

//BADD_2397 replaced by BADD_2820

//BADD_2396 replaced by BADD_2819

//BADD_2395 replaced by BADD_2818

//ADD_7386 replaced by ADD_8288

//ADD_7385 replaced by ADD_8288

//KaratsubaCore_1079 replaced by KaratsubaCore_1438

//KaratsubaCore_1078 replaced by KaratsubaCore_1435

//KaratsubaCore_1077 replaced by KaratsubaCore_1438

//ADD_7392 replaced by ADD_11602

//ADD_7391 replaced by ADD_11602

//ADD_7390 replaced by ADD_11602

//ADD_7389 replaced by ADD_11602

//ADD_7388 replaced by ADD_11602

//ADD_7387 replaced by ADD_11602

//ADD_7397 replaced by ADD_11601

//ADD_7396 replaced by ADD_11602

//ADD_7395 replaced by ADD_11602

//ADD_7394 replaced by ADD_11602

//ADD_7393 replaced by ADD_11602

//ADD_7401 replaced by ADD_11602

//ADD_7400 replaced by ADD_11602

//ADD_7399 replaced by ADD_11602

//ADD_7398 replaced by ADD_11602

//BADD_2401 replaced by BADD_2824

//BADD_2400 replaced by BADD_2823

//BADD_2399 replaced by BADD_2822

//ADD_7403 replaced by ADD_11602

//ADD_7402 replaced by ADD_11602

//KaratsubaCore_1082 replaced by KaratsubaCore_1437

//KaratsubaCore_1081 replaced by KaratsubaCore_1438

//KaratsubaCore_1080 replaced by KaratsubaCore_1437

//BADD_2405 replaced by BADD_2818

//BADD_2404 replaced by BADD_2820

//BADD_2403 replaced by BADD_2819

//BADD_2402 replaced by BADD_2818

//ADD_7405 replaced by ADD_8288

//ADD_7404 replaced by ADD_8288

//KaratsubaCore_1085 replaced by KaratsubaCore_1438

//KaratsubaCore_1084 replaced by KaratsubaCore_1435

//KaratsubaCore_1083 replaced by KaratsubaCore_1438

//BADD_2408 replaced by BADD_2824

//BADD_2407 replaced by BADD_2823

//BADD_2406 replaced by BADD_2822

//ADD_7407 replaced by ADD_11602

//ADD_7406 replaced by ADD_11602

//KaratsubaCore_1088 replaced by KaratsubaCore_1437

//KaratsubaCore_1087 replaced by KaratsubaCore_1438

//KaratsubaCore_1086 replaced by KaratsubaCore_1437

//ADD_7413 replaced by ADD_11602

//ADD_7412 replaced by ADD_11602

//ADD_7411 replaced by ADD_11602

//ADD_7410 replaced by ADD_11602

//ADD_7409 replaced by ADD_11602

//ADD_7408 replaced by ADD_11602

//ADD_7418 replaced by ADD_11601

//ADD_7417 replaced by ADD_11602

//ADD_7416 replaced by ADD_11602

//ADD_7415 replaced by ADD_11602

//ADD_7414 replaced by ADD_11602

//ADD_7422 replaced by ADD_11602

//ADD_7421 replaced by ADD_11602

//ADD_7420 replaced by ADD_11602

//ADD_7419 replaced by ADD_11602

//BADD_2411 replaced by BADD_2824

//BADD_2410 replaced by BADD_2823

//BADD_2409 replaced by BADD_2822

//ADD_7424 replaced by ADD_11602

//ADD_7423 replaced by ADD_11602

//KaratsubaCore_1091 replaced by KaratsubaCore_1437

//KaratsubaCore_1090 replaced by KaratsubaCore_1438

//KaratsubaCore_1089 replaced by KaratsubaCore_1437

//BADD_2415 replaced by BADD_2818

//BADD_2414 replaced by BADD_2820

//BADD_2413 replaced by BADD_2819

//BADD_2412 replaced by BADD_2818

//ADD_7426 replaced by ADD_8288

//ADD_7425 replaced by ADD_8288

//KaratsubaCore_1094 replaced by KaratsubaCore_1438

//KaratsubaCore_1093 replaced by KaratsubaCore_1435

//KaratsubaCore_1092 replaced by KaratsubaCore_1438

//BADD_2418 replaced by BADD_2824

//BADD_2417 replaced by BADD_2823

//BADD_2416 replaced by BADD_2822

//ADD_7428 replaced by ADD_11602

//ADD_7427 replaced by ADD_11602

//KaratsubaCore_1097 replaced by KaratsubaCore_1437

//KaratsubaCore_1096 replaced by KaratsubaCore_1438

//KaratsubaCore_1095 replaced by KaratsubaCore_1437

//ADD_7433 replaced by ADD_11595

//ADD_7432 replaced by ADD_11602

//ADD_7431 replaced by ADD_11602

//ADD_7430 replaced by ADD_11602

//ADD_7429 replaced by ADD_11602

//ADD_7438 replaced by ADD_11592

//ADD_7437 replaced by ADD_11602

//ADD_7436 replaced by ADD_11602

//ADD_7435 replaced by ADD_11602

//ADD_7434 replaced by ADD_11602

//ADD_7443 replaced by ADD_11592

//ADD_7442 replaced by ADD_11602

//ADD_7441 replaced by ADD_11602

//ADD_7440 replaced by ADD_11602

//ADD_7439 replaced by ADD_11602

//ADD_7448 replaced by ADD_11595

//ADD_7447 replaced by ADD_11602

//ADD_7446 replaced by ADD_11602

//ADD_7445 replaced by ADD_11602

//ADD_7444 replaced by ADD_11602

//BADD_2422 replaced by BADD_2818

//BADD_2421 replaced by BADD_2820

//BADD_2420 replaced by BADD_2819

//BADD_2419 replaced by BADD_2818

//ADD_7450 replaced by ADD_8288

//ADD_7449 replaced by ADD_8288

//KaratsubaCore_1100 replaced by KaratsubaCore_1438

//KaratsubaCore_1099 replaced by KaratsubaCore_1435

//KaratsubaCore_1098 replaced by KaratsubaCore_1438

//BADD_2426 replaced by BADD_2807

//BADD_2425 replaced by BADD_2809

//BADD_2424 replaced by BADD_2808

//BADD_2423 replaced by BADD_2807

//ADD_7452 replaced by ADD_8267

//ADD_7451 replaced by ADD_8267

//KaratsubaCore_1103 replaced by KaratsubaCore_1435

//KaratsubaCore_1102 replaced by KaratsubaCore_1426

//KaratsubaCore_1101 replaced by KaratsubaCore_1435

//BADD_2430 replaced by BADD_2818

//BADD_2429 replaced by BADD_2820

//BADD_2428 replaced by BADD_2819

//BADD_2427 replaced by BADD_2818

//ADD_7454 replaced by ADD_8288

//ADD_7453 replaced by ADD_8288

//KaratsubaCore_1106 replaced by KaratsubaCore_1438

//KaratsubaCore_1105 replaced by KaratsubaCore_1435

//KaratsubaCore_1104 replaced by KaratsubaCore_1438

//ADD_7460 replaced by ADD_11602

//ADD_7459 replaced by ADD_11602

//ADD_7458 replaced by ADD_11602

//ADD_7457 replaced by ADD_11602

//ADD_7456 replaced by ADD_11602

//ADD_7455 replaced by ADD_11602

//ADD_7465 replaced by ADD_11601

//ADD_7464 replaced by ADD_11602

//ADD_7463 replaced by ADD_11602

//ADD_7462 replaced by ADD_11602

//ADD_7461 replaced by ADD_11602

//ADD_7469 replaced by ADD_11602

//ADD_7468 replaced by ADD_11602

//ADD_7467 replaced by ADD_11602

//ADD_7466 replaced by ADD_11602

//BADD_2433 replaced by BADD_2824

//BADD_2432 replaced by BADD_2823

//BADD_2431 replaced by BADD_2822

//ADD_7471 replaced by ADD_11602

//ADD_7470 replaced by ADD_11602

//KaratsubaCore_1109 replaced by KaratsubaCore_1437

//KaratsubaCore_1108 replaced by KaratsubaCore_1438

//KaratsubaCore_1107 replaced by KaratsubaCore_1437

//BADD_2437 replaced by BADD_2818

//BADD_2436 replaced by BADD_2820

//BADD_2435 replaced by BADD_2819

//BADD_2434 replaced by BADD_2818

//ADD_7473 replaced by ADD_8288

//ADD_7472 replaced by ADD_8288

//KaratsubaCore_1112 replaced by KaratsubaCore_1438

//KaratsubaCore_1111 replaced by KaratsubaCore_1435

//KaratsubaCore_1110 replaced by KaratsubaCore_1438

//BADD_2440 replaced by BADD_2824

//BADD_2439 replaced by BADD_2823

//BADD_2438 replaced by BADD_2822

//ADD_7475 replaced by ADD_11602

//ADD_7474 replaced by ADD_11602

//KaratsubaCore_1115 replaced by KaratsubaCore_1437

//KaratsubaCore_1114 replaced by KaratsubaCore_1438

//KaratsubaCore_1113 replaced by KaratsubaCore_1437

//ADD_7481 replaced by ADD_11602

//ADD_7480 replaced by ADD_11602

//ADD_7479 replaced by ADD_11602

//ADD_7478 replaced by ADD_11602

//ADD_7477 replaced by ADD_11602

//ADD_7476 replaced by ADD_11602

//ADD_7486 replaced by ADD_11601

//ADD_7485 replaced by ADD_11602

//ADD_7484 replaced by ADD_11602

//ADD_7483 replaced by ADD_11602

//ADD_7482 replaced by ADD_11602

//ADD_7490 replaced by ADD_11602

//ADD_7489 replaced by ADD_11602

//ADD_7488 replaced by ADD_11602

//ADD_7487 replaced by ADD_11602

//BADD_2443 replaced by BADD_2824

//BADD_2442 replaced by BADD_2823

//BADD_2441 replaced by BADD_2822

//ADD_7492 replaced by ADD_11602

//ADD_7491 replaced by ADD_11602

//KaratsubaCore_1118 replaced by KaratsubaCore_1437

//KaratsubaCore_1117 replaced by KaratsubaCore_1438

//KaratsubaCore_1116 replaced by KaratsubaCore_1437

//BADD_2447 replaced by BADD_2818

//BADD_2446 replaced by BADD_2820

//BADD_2445 replaced by BADD_2819

//BADD_2444 replaced by BADD_2818

//ADD_7494 replaced by ADD_8288

//ADD_7493 replaced by ADD_8288

//KaratsubaCore_1121 replaced by KaratsubaCore_1438

//KaratsubaCore_1120 replaced by KaratsubaCore_1435

//KaratsubaCore_1119 replaced by KaratsubaCore_1438

//BADD_2450 replaced by BADD_2824

//BADD_2449 replaced by BADD_2823

//BADD_2448 replaced by BADD_2822

//ADD_7496 replaced by ADD_11602

//ADD_7495 replaced by ADD_11602

//KaratsubaCore_1124 replaced by KaratsubaCore_1437

//KaratsubaCore_1123 replaced by KaratsubaCore_1438

//KaratsubaCore_1122 replaced by KaratsubaCore_1437

//ADD_7501 replaced by ADD_11595

//ADD_7500 replaced by ADD_11602

//ADD_7499 replaced by ADD_11602

//ADD_7498 replaced by ADD_11602

//ADD_7497 replaced by ADD_11602

//ADD_7506 replaced by ADD_11592

//ADD_7505 replaced by ADD_11602

//ADD_7504 replaced by ADD_11602

//ADD_7503 replaced by ADD_11602

//ADD_7502 replaced by ADD_11602

//ADD_7511 replaced by ADD_11592

//ADD_7510 replaced by ADD_11602

//ADD_7509 replaced by ADD_11602

//ADD_7508 replaced by ADD_11602

//ADD_7507 replaced by ADD_11602

//ADD_7516 replaced by ADD_11595

//ADD_7515 replaced by ADD_11602

//ADD_7514 replaced by ADD_11602

//ADD_7513 replaced by ADD_11602

//ADD_7512 replaced by ADD_11602

//BADD_2454 replaced by BADD_2818

//BADD_2453 replaced by BADD_2820

//BADD_2452 replaced by BADD_2819

//BADD_2451 replaced by BADD_2818

//ADD_7518 replaced by ADD_8288

//ADD_7517 replaced by ADD_8288

//KaratsubaCore_1127 replaced by KaratsubaCore_1438

//KaratsubaCore_1126 replaced by KaratsubaCore_1435

//KaratsubaCore_1125 replaced by KaratsubaCore_1438

//BADD_2458 replaced by BADD_2807

//BADD_2457 replaced by BADD_2809

//BADD_2456 replaced by BADD_2808

//BADD_2455 replaced by BADD_2807

//ADD_7520 replaced by ADD_8267

//ADD_7519 replaced by ADD_8267

//KaratsubaCore_1130 replaced by KaratsubaCore_1435

//KaratsubaCore_1129 replaced by KaratsubaCore_1426

//KaratsubaCore_1128 replaced by KaratsubaCore_1435

//BADD_2462 replaced by BADD_2818

//BADD_2461 replaced by BADD_2820

//BADD_2460 replaced by BADD_2819

//BADD_2459 replaced by BADD_2818

//ADD_7522 replaced by ADD_8288

//ADD_7521 replaced by ADD_8288

//KaratsubaCore_1133 replaced by KaratsubaCore_1438

//KaratsubaCore_1132 replaced by KaratsubaCore_1435

//KaratsubaCore_1131 replaced by KaratsubaCore_1438

//ADD_7528 replaced by ADD_11602

//ADD_7527 replaced by ADD_11602

//ADD_7526 replaced by ADD_11602

//ADD_7525 replaced by ADD_11602

//ADD_7524 replaced by ADD_11602

//ADD_7523 replaced by ADD_11602

//ADD_7533 replaced by ADD_11601

//ADD_7532 replaced by ADD_11602

//ADD_7531 replaced by ADD_11602

//ADD_7530 replaced by ADD_11602

//ADD_7529 replaced by ADD_11602

//ADD_7537 replaced by ADD_11602

//ADD_7536 replaced by ADD_11602

//ADD_7535 replaced by ADD_11602

//ADD_7534 replaced by ADD_11602

//BADD_2465 replaced by BADD_2824

//BADD_2464 replaced by BADD_2823

//BADD_2463 replaced by BADD_2822

//ADD_7539 replaced by ADD_11602

//ADD_7538 replaced by ADD_11602

//KaratsubaCore_1136 replaced by KaratsubaCore_1437

//KaratsubaCore_1135 replaced by KaratsubaCore_1438

//KaratsubaCore_1134 replaced by KaratsubaCore_1437

//BADD_2469 replaced by BADD_2818

//BADD_2468 replaced by BADD_2820

//BADD_2467 replaced by BADD_2819

//BADD_2466 replaced by BADD_2818

//ADD_7541 replaced by ADD_8288

//ADD_7540 replaced by ADD_8288

//KaratsubaCore_1139 replaced by KaratsubaCore_1438

//KaratsubaCore_1138 replaced by KaratsubaCore_1435

//KaratsubaCore_1137 replaced by KaratsubaCore_1438

//BADD_2472 replaced by BADD_2824

//BADD_2471 replaced by BADD_2823

//BADD_2470 replaced by BADD_2822

//ADD_7543 replaced by ADD_11602

//ADD_7542 replaced by ADD_11602

//KaratsubaCore_1142 replaced by KaratsubaCore_1437

//KaratsubaCore_1141 replaced by KaratsubaCore_1438

//KaratsubaCore_1140 replaced by KaratsubaCore_1437

//ADD_7549 replaced by ADD_11602

//ADD_7548 replaced by ADD_11602

//ADD_7547 replaced by ADD_11602

//ADD_7546 replaced by ADD_11602

//ADD_7545 replaced by ADD_11602

//ADD_7544 replaced by ADD_11602

//ADD_7554 replaced by ADD_11601

//ADD_7553 replaced by ADD_11602

//ADD_7552 replaced by ADD_11602

//ADD_7551 replaced by ADD_11602

//ADD_7550 replaced by ADD_11602

//ADD_7558 replaced by ADD_11602

//ADD_7557 replaced by ADD_11602

//ADD_7556 replaced by ADD_11602

//ADD_7555 replaced by ADD_11602

//BADD_2475 replaced by BADD_2824

//BADD_2474 replaced by BADD_2823

//BADD_2473 replaced by BADD_2822

//ADD_7560 replaced by ADD_11602

//ADD_7559 replaced by ADD_11602

//KaratsubaCore_1145 replaced by KaratsubaCore_1437

//KaratsubaCore_1144 replaced by KaratsubaCore_1438

//KaratsubaCore_1143 replaced by KaratsubaCore_1437

//BADD_2479 replaced by BADD_2818

//BADD_2478 replaced by BADD_2820

//BADD_2477 replaced by BADD_2819

//BADD_2476 replaced by BADD_2818

//ADD_7562 replaced by ADD_8288

//ADD_7561 replaced by ADD_8288

//KaratsubaCore_1148 replaced by KaratsubaCore_1438

//KaratsubaCore_1147 replaced by KaratsubaCore_1435

//KaratsubaCore_1146 replaced by KaratsubaCore_1438

//BADD_2482 replaced by BADD_2824

//BADD_2481 replaced by BADD_2823

//BADD_2480 replaced by BADD_2822

//ADD_7564 replaced by ADD_11602

//ADD_7563 replaced by ADD_11602

//KaratsubaCore_1151 replaced by KaratsubaCore_1437

//KaratsubaCore_1150 replaced by KaratsubaCore_1438

//KaratsubaCore_1149 replaced by KaratsubaCore_1437

//ADD_7569 replaced by ADD_11595

//ADD_7568 replaced by ADD_11602

//ADD_7567 replaced by ADD_11602

//ADD_7566 replaced by ADD_11602

//ADD_7565 replaced by ADD_11602

//ADD_7574 replaced by ADD_11592

//ADD_7573 replaced by ADD_11602

//ADD_7572 replaced by ADD_11602

//ADD_7571 replaced by ADD_11602

//ADD_7570 replaced by ADD_11602

//ADD_7579 replaced by ADD_11592

//ADD_7578 replaced by ADD_11602

//ADD_7577 replaced by ADD_11602

//ADD_7576 replaced by ADD_11602

//ADD_7575 replaced by ADD_11602

//ADD_7584 replaced by ADD_11595

//ADD_7583 replaced by ADD_11602

//ADD_7582 replaced by ADD_11602

//ADD_7581 replaced by ADD_11602

//ADD_7580 replaced by ADD_11602

//BADD_2486 replaced by BADD_2818

//BADD_2485 replaced by BADD_2820

//BADD_2484 replaced by BADD_2819

//BADD_2483 replaced by BADD_2818

//ADD_7586 replaced by ADD_8288

//ADD_7585 replaced by ADD_8288

//KaratsubaCore_1154 replaced by KaratsubaCore_1438

//KaratsubaCore_1153 replaced by KaratsubaCore_1435

//KaratsubaCore_1152 replaced by KaratsubaCore_1438

//BADD_2490 replaced by BADD_2807

//BADD_2489 replaced by BADD_2809

//BADD_2488 replaced by BADD_2808

//BADD_2487 replaced by BADD_2807

//ADD_7588 replaced by ADD_8267

//ADD_7587 replaced by ADD_8267

//KaratsubaCore_1157 replaced by KaratsubaCore_1435

//KaratsubaCore_1156 replaced by KaratsubaCore_1426

//KaratsubaCore_1155 replaced by KaratsubaCore_1435

//BADD_2494 replaced by BADD_2818

//BADD_2493 replaced by BADD_2820

//BADD_2492 replaced by BADD_2819

//BADD_2491 replaced by BADD_2818

//ADD_7590 replaced by ADD_8288

//ADD_7589 replaced by ADD_8288

//KaratsubaCore_1160 replaced by KaratsubaCore_1438

//KaratsubaCore_1159 replaced by KaratsubaCore_1435

//KaratsubaCore_1158 replaced by KaratsubaCore_1438

//ADD_7596 replaced by ADD_11602

//ADD_7595 replaced by ADD_11602

//ADD_7594 replaced by ADD_11602

//ADD_7593 replaced by ADD_11602

//ADD_7592 replaced by ADD_11602

//ADD_7591 replaced by ADD_11602

//ADD_7601 replaced by ADD_11601

//ADD_7600 replaced by ADD_11602

//ADD_7599 replaced by ADD_11602

//ADD_7598 replaced by ADD_11602

//ADD_7597 replaced by ADD_11602

//ADD_7605 replaced by ADD_11602

//ADD_7604 replaced by ADD_11602

//ADD_7603 replaced by ADD_11602

//ADD_7602 replaced by ADD_11602

//BADD_2497 replaced by BADD_2824

//BADD_2496 replaced by BADD_2823

//BADD_2495 replaced by BADD_2822

//ADD_7607 replaced by ADD_11602

//ADD_7606 replaced by ADD_11602

//KaratsubaCore_1163 replaced by KaratsubaCore_1437

//KaratsubaCore_1162 replaced by KaratsubaCore_1438

//KaratsubaCore_1161 replaced by KaratsubaCore_1437

//BADD_2501 replaced by BADD_2818

//BADD_2500 replaced by BADD_2820

//BADD_2499 replaced by BADD_2819

//BADD_2498 replaced by BADD_2818

//ADD_7609 replaced by ADD_8288

//ADD_7608 replaced by ADD_8288

//KaratsubaCore_1166 replaced by KaratsubaCore_1438

//KaratsubaCore_1165 replaced by KaratsubaCore_1435

//KaratsubaCore_1164 replaced by KaratsubaCore_1438

//BADD_2504 replaced by BADD_2824

//BADD_2503 replaced by BADD_2823

//BADD_2502 replaced by BADD_2822

//ADD_7611 replaced by ADD_11602

//ADD_7610 replaced by ADD_11602

//KaratsubaCore_1169 replaced by KaratsubaCore_1437

//KaratsubaCore_1168 replaced by KaratsubaCore_1438

//KaratsubaCore_1167 replaced by KaratsubaCore_1437

//ADD_7617 replaced by ADD_11602

//ADD_7616 replaced by ADD_11602

//ADD_7615 replaced by ADD_11602

//ADD_7614 replaced by ADD_11602

//ADD_7613 replaced by ADD_11602

//ADD_7612 replaced by ADD_11602

//ADD_7622 replaced by ADD_11601

//ADD_7621 replaced by ADD_11602

//ADD_7620 replaced by ADD_11602

//ADD_7619 replaced by ADD_11602

//ADD_7618 replaced by ADD_11602

//ADD_7626 replaced by ADD_11602

//ADD_7625 replaced by ADD_11602

//ADD_7624 replaced by ADD_11602

//ADD_7623 replaced by ADD_11602

//BADD_2507 replaced by BADD_2824

//BADD_2506 replaced by BADD_2823

//BADD_2505 replaced by BADD_2822

//ADD_7628 replaced by ADD_11602

//ADD_7627 replaced by ADD_11602

//KaratsubaCore_1172 replaced by KaratsubaCore_1437

//KaratsubaCore_1171 replaced by KaratsubaCore_1438

//KaratsubaCore_1170 replaced by KaratsubaCore_1437

//BADD_2511 replaced by BADD_2818

//BADD_2510 replaced by BADD_2820

//BADD_2509 replaced by BADD_2819

//BADD_2508 replaced by BADD_2818

//ADD_7630 replaced by ADD_8288

//ADD_7629 replaced by ADD_8288

//KaratsubaCore_1175 replaced by KaratsubaCore_1438

//KaratsubaCore_1174 replaced by KaratsubaCore_1435

//KaratsubaCore_1173 replaced by KaratsubaCore_1438

//BADD_2514 replaced by BADD_2824

//BADD_2513 replaced by BADD_2823

//BADD_2512 replaced by BADD_2822

//ADD_7632 replaced by ADD_11602

//ADD_7631 replaced by ADD_11602

//KaratsubaCore_1178 replaced by KaratsubaCore_1437

//KaratsubaCore_1177 replaced by KaratsubaCore_1438

//KaratsubaCore_1176 replaced by KaratsubaCore_1437

//ADD_7637 replaced by ADD_11595

//ADD_7636 replaced by ADD_11602

//ADD_7635 replaced by ADD_11602

//ADD_7634 replaced by ADD_11602

//ADD_7633 replaced by ADD_11602

//ADD_7642 replaced by ADD_11592

//ADD_7641 replaced by ADD_11602

//ADD_7640 replaced by ADD_11602

//ADD_7639 replaced by ADD_11602

//ADD_7638 replaced by ADD_11602

//ADD_7647 replaced by ADD_11592

//ADD_7646 replaced by ADD_11602

//ADD_7645 replaced by ADD_11602

//ADD_7644 replaced by ADD_11602

//ADD_7643 replaced by ADD_11602

//ADD_7652 replaced by ADD_11595

//ADD_7651 replaced by ADD_11602

//ADD_7650 replaced by ADD_11602

//ADD_7649 replaced by ADD_11602

//ADD_7648 replaced by ADD_11602

//BADD_2518 replaced by BADD_2818

//BADD_2517 replaced by BADD_2820

//BADD_2516 replaced by BADD_2819

//BADD_2515 replaced by BADD_2818

//ADD_7654 replaced by ADD_8288

//ADD_7653 replaced by ADD_8288

//KaratsubaCore_1181 replaced by KaratsubaCore_1438

//KaratsubaCore_1180 replaced by KaratsubaCore_1435

//KaratsubaCore_1179 replaced by KaratsubaCore_1438

//BADD_2522 replaced by BADD_2807

//BADD_2521 replaced by BADD_2809

//BADD_2520 replaced by BADD_2808

//BADD_2519 replaced by BADD_2807

//ADD_7656 replaced by ADD_8267

//ADD_7655 replaced by ADD_8267

//KaratsubaCore_1184 replaced by KaratsubaCore_1435

//KaratsubaCore_1183 replaced by KaratsubaCore_1426

//KaratsubaCore_1182 replaced by KaratsubaCore_1435

//BADD_2526 replaced by BADD_2818

//BADD_2525 replaced by BADD_2820

//BADD_2524 replaced by BADD_2819

//BADD_2523 replaced by BADD_2818

//ADD_7658 replaced by ADD_8288

//ADD_7657 replaced by ADD_8288

//KaratsubaCore_1187 replaced by KaratsubaCore_1438

//KaratsubaCore_1186 replaced by KaratsubaCore_1435

//KaratsubaCore_1185 replaced by KaratsubaCore_1438

//ADD_7664 replaced by ADD_11602

//ADD_7663 replaced by ADD_11602

//ADD_7662 replaced by ADD_11602

//ADD_7661 replaced by ADD_11602

//ADD_7660 replaced by ADD_11602

//ADD_7659 replaced by ADD_11602

//ADD_7669 replaced by ADD_11601

//ADD_7668 replaced by ADD_11602

//ADD_7667 replaced by ADD_11602

//ADD_7666 replaced by ADD_11602

//ADD_7665 replaced by ADD_11602

//ADD_7673 replaced by ADD_11602

//ADD_7672 replaced by ADD_11602

//ADD_7671 replaced by ADD_11602

//ADD_7670 replaced by ADD_11602

//BADD_2529 replaced by BADD_2824

//BADD_2528 replaced by BADD_2823

//BADD_2527 replaced by BADD_2822

//ADD_7675 replaced by ADD_11602

//ADD_7674 replaced by ADD_11602

//KaratsubaCore_1190 replaced by KaratsubaCore_1437

//KaratsubaCore_1189 replaced by KaratsubaCore_1438

//KaratsubaCore_1188 replaced by KaratsubaCore_1437

//BADD_2533 replaced by BADD_2818

//BADD_2532 replaced by BADD_2820

//BADD_2531 replaced by BADD_2819

//BADD_2530 replaced by BADD_2818

//ADD_7677 replaced by ADD_8288

//ADD_7676 replaced by ADD_8288

//KaratsubaCore_1193 replaced by KaratsubaCore_1438

//KaratsubaCore_1192 replaced by KaratsubaCore_1435

//KaratsubaCore_1191 replaced by KaratsubaCore_1438

//BADD_2536 replaced by BADD_2824

//BADD_2535 replaced by BADD_2823

//BADD_2534 replaced by BADD_2822

//ADD_7679 replaced by ADD_11602

//ADD_7678 replaced by ADD_11602

//KaratsubaCore_1196 replaced by KaratsubaCore_1437

//KaratsubaCore_1195 replaced by KaratsubaCore_1438

//KaratsubaCore_1194 replaced by KaratsubaCore_1437

//ADD_7685 replaced by ADD_11602

//ADD_7684 replaced by ADD_11602

//ADD_7683 replaced by ADD_11602

//ADD_7682 replaced by ADD_11602

//ADD_7681 replaced by ADD_11602

//ADD_7680 replaced by ADD_11602

//ADD_7690 replaced by ADD_11601

//ADD_7689 replaced by ADD_11602

//ADD_7688 replaced by ADD_11602

//ADD_7687 replaced by ADD_11602

//ADD_7686 replaced by ADD_11602

//ADD_7694 replaced by ADD_11602

//ADD_7693 replaced by ADD_11602

//ADD_7692 replaced by ADD_11602

//ADD_7691 replaced by ADD_11602

//BADD_2539 replaced by BADD_2824

//BADD_2538 replaced by BADD_2823

//BADD_2537 replaced by BADD_2822

//ADD_7696 replaced by ADD_11602

//ADD_7695 replaced by ADD_11602

//KaratsubaCore_1199 replaced by KaratsubaCore_1437

//KaratsubaCore_1198 replaced by KaratsubaCore_1438

//KaratsubaCore_1197 replaced by KaratsubaCore_1437

//BADD_2543 replaced by BADD_2818

//BADD_2542 replaced by BADD_2820

//BADD_2541 replaced by BADD_2819

//BADD_2540 replaced by BADD_2818

//ADD_7698 replaced by ADD_8288

//ADD_7697 replaced by ADD_8288

//KaratsubaCore_1202 replaced by KaratsubaCore_1438

//KaratsubaCore_1201 replaced by KaratsubaCore_1435

//KaratsubaCore_1200 replaced by KaratsubaCore_1438

//BADD_2546 replaced by BADD_2824

//BADD_2545 replaced by BADD_2823

//BADD_2544 replaced by BADD_2822

//ADD_7700 replaced by ADD_11602

//ADD_7699 replaced by ADD_11602

//KaratsubaCore_1205 replaced by KaratsubaCore_1437

//KaratsubaCore_1204 replaced by KaratsubaCore_1438

//KaratsubaCore_1203 replaced by KaratsubaCore_1437

//ADD_7705 replaced by ADD_11595

//ADD_7704 replaced by ADD_11602

//ADD_7703 replaced by ADD_11602

//ADD_7702 replaced by ADD_11602

//ADD_7701 replaced by ADD_11602

//ADD_7710 replaced by ADD_11592

//ADD_7709 replaced by ADD_11602

//ADD_7708 replaced by ADD_11602

//ADD_7707 replaced by ADD_11602

//ADD_7706 replaced by ADD_11602

//ADD_7715 replaced by ADD_11592

//ADD_7714 replaced by ADD_11602

//ADD_7713 replaced by ADD_11602

//ADD_7712 replaced by ADD_11602

//ADD_7711 replaced by ADD_11602

//ADD_7720 replaced by ADD_11595

//ADD_7719 replaced by ADD_11602

//ADD_7718 replaced by ADD_11602

//ADD_7717 replaced by ADD_11602

//ADD_7716 replaced by ADD_11602

//BADD_2550 replaced by BADD_2818

//BADD_2549 replaced by BADD_2820

//BADD_2548 replaced by BADD_2819

//BADD_2547 replaced by BADD_2818

//ADD_7722 replaced by ADD_8288

//ADD_7721 replaced by ADD_8288

//KaratsubaCore_1208 replaced by KaratsubaCore_1438

//KaratsubaCore_1207 replaced by KaratsubaCore_1435

//KaratsubaCore_1206 replaced by KaratsubaCore_1438

//BADD_2554 replaced by BADD_2807

//BADD_2553 replaced by BADD_2809

//BADD_2552 replaced by BADD_2808

//BADD_2551 replaced by BADD_2807

//ADD_7724 replaced by ADD_8267

//ADD_7723 replaced by ADD_8267

//KaratsubaCore_1211 replaced by KaratsubaCore_1435

//KaratsubaCore_1210 replaced by KaratsubaCore_1426

//KaratsubaCore_1209 replaced by KaratsubaCore_1435

//BADD_2558 replaced by BADD_2818

//BADD_2557 replaced by BADD_2820

//BADD_2556 replaced by BADD_2819

//BADD_2555 replaced by BADD_2818

//ADD_7726 replaced by ADD_8288

//ADD_7725 replaced by ADD_8288

//KaratsubaCore_1214 replaced by KaratsubaCore_1438

//KaratsubaCore_1213 replaced by KaratsubaCore_1435

//KaratsubaCore_1212 replaced by KaratsubaCore_1438

//ADD_7732 replaced by ADD_11602

//ADD_7731 replaced by ADD_11602

//ADD_7730 replaced by ADD_11602

//ADD_7729 replaced by ADD_11602

//ADD_7728 replaced by ADD_11602

//ADD_7727 replaced by ADD_11602

//ADD_7737 replaced by ADD_11601

//ADD_7736 replaced by ADD_11602

//ADD_7735 replaced by ADD_11602

//ADD_7734 replaced by ADD_11602

//ADD_7733 replaced by ADD_11602

//ADD_7741 replaced by ADD_11602

//ADD_7740 replaced by ADD_11602

//ADD_7739 replaced by ADD_11602

//ADD_7738 replaced by ADD_11602

//BADD_2561 replaced by BADD_2824

//BADD_2560 replaced by BADD_2823

//BADD_2559 replaced by BADD_2822

//ADD_7743 replaced by ADD_11602

//ADD_7742 replaced by ADD_11602

//KaratsubaCore_1217 replaced by KaratsubaCore_1437

//KaratsubaCore_1216 replaced by KaratsubaCore_1438

//KaratsubaCore_1215 replaced by KaratsubaCore_1437

//BADD_2565 replaced by BADD_2818

//BADD_2564 replaced by BADD_2820

//BADD_2563 replaced by BADD_2819

//BADD_2562 replaced by BADD_2818

//ADD_7745 replaced by ADD_8288

//ADD_7744 replaced by ADD_8288

//KaratsubaCore_1220 replaced by KaratsubaCore_1438

//KaratsubaCore_1219 replaced by KaratsubaCore_1435

//KaratsubaCore_1218 replaced by KaratsubaCore_1438

//BADD_2568 replaced by BADD_2824

//BADD_2567 replaced by BADD_2823

//BADD_2566 replaced by BADD_2822

//ADD_7747 replaced by ADD_11602

//ADD_7746 replaced by ADD_11602

//KaratsubaCore_1223 replaced by KaratsubaCore_1437

//KaratsubaCore_1222 replaced by KaratsubaCore_1438

//KaratsubaCore_1221 replaced by KaratsubaCore_1437

//ADD_7753 replaced by ADD_11602

//ADD_7752 replaced by ADD_11602

//ADD_7751 replaced by ADD_11602

//ADD_7750 replaced by ADD_11602

//ADD_7749 replaced by ADD_11602

//ADD_7748 replaced by ADD_11602

//ADD_7758 replaced by ADD_11601

//ADD_7757 replaced by ADD_11602

//ADD_7756 replaced by ADD_11602

//ADD_7755 replaced by ADD_11602

//ADD_7754 replaced by ADD_11602

//ADD_7762 replaced by ADD_11602

//ADD_7761 replaced by ADD_11602

//ADD_7760 replaced by ADD_11602

//ADD_7759 replaced by ADD_11602

//BADD_2571 replaced by BADD_2824

//BADD_2570 replaced by BADD_2823

//BADD_2569 replaced by BADD_2822

//ADD_7764 replaced by ADD_11602

//ADD_7763 replaced by ADD_11602

//KaratsubaCore_1226 replaced by KaratsubaCore_1437

//KaratsubaCore_1225 replaced by KaratsubaCore_1438

//KaratsubaCore_1224 replaced by KaratsubaCore_1437

//BADD_2575 replaced by BADD_2818

//BADD_2574 replaced by BADD_2820

//BADD_2573 replaced by BADD_2819

//BADD_2572 replaced by BADD_2818

//ADD_7766 replaced by ADD_8288

//ADD_7765 replaced by ADD_8288

//KaratsubaCore_1229 replaced by KaratsubaCore_1438

//KaratsubaCore_1228 replaced by KaratsubaCore_1435

//KaratsubaCore_1227 replaced by KaratsubaCore_1438

//BADD_2578 replaced by BADD_2824

//BADD_2577 replaced by BADD_2823

//BADD_2576 replaced by BADD_2822

//ADD_7768 replaced by ADD_11602

//ADD_7767 replaced by ADD_11602

//KaratsubaCore_1232 replaced by KaratsubaCore_1437

//KaratsubaCore_1231 replaced by KaratsubaCore_1438

//KaratsubaCore_1230 replaced by KaratsubaCore_1437

//ADD_7773 replaced by ADD_11595

//ADD_7772 replaced by ADD_11602

//ADD_7771 replaced by ADD_11602

//ADD_7770 replaced by ADD_11602

//ADD_7769 replaced by ADD_11602

//ADD_7778 replaced by ADD_11592

//ADD_7777 replaced by ADD_11602

//ADD_7776 replaced by ADD_11602

//ADD_7775 replaced by ADD_11602

//ADD_7774 replaced by ADD_11602

//ADD_7783 replaced by ADD_11592

//ADD_7782 replaced by ADD_11602

//ADD_7781 replaced by ADD_11602

//ADD_7780 replaced by ADD_11602

//ADD_7779 replaced by ADD_11602

//ADD_7788 replaced by ADD_11595

//ADD_7787 replaced by ADD_11602

//ADD_7786 replaced by ADD_11602

//ADD_7785 replaced by ADD_11602

//ADD_7784 replaced by ADD_11602

//BADD_2582 replaced by BADD_2818

//BADD_2581 replaced by BADD_2820

//BADD_2580 replaced by BADD_2819

//BADD_2579 replaced by BADD_2818

//ADD_7790 replaced by ADD_8288

//ADD_7789 replaced by ADD_8288

//KaratsubaCore_1235 replaced by KaratsubaCore_1438

//KaratsubaCore_1234 replaced by KaratsubaCore_1435

//KaratsubaCore_1233 replaced by KaratsubaCore_1438

//BADD_2586 replaced by BADD_2807

//BADD_2585 replaced by BADD_2809

//BADD_2584 replaced by BADD_2808

//BADD_2583 replaced by BADD_2807

//ADD_7792 replaced by ADD_8267

//ADD_7791 replaced by ADD_8267

//KaratsubaCore_1238 replaced by KaratsubaCore_1435

//KaratsubaCore_1237 replaced by KaratsubaCore_1426

//KaratsubaCore_1236 replaced by KaratsubaCore_1435

//BADD_2590 replaced by BADD_2818

//BADD_2589 replaced by BADD_2820

//BADD_2588 replaced by BADD_2819

//BADD_2587 replaced by BADD_2818

//ADD_7794 replaced by ADD_8288

//ADD_7793 replaced by ADD_8288

//KaratsubaCore_1241 replaced by KaratsubaCore_1438

//KaratsubaCore_1240 replaced by KaratsubaCore_1435

//KaratsubaCore_1239 replaced by KaratsubaCore_1438

//ADD_7800 replaced by ADD_11602

//ADD_7799 replaced by ADD_11602

//ADD_7798 replaced by ADD_11602

//ADD_7797 replaced by ADD_11602

//ADD_7796 replaced by ADD_11602

//ADD_7795 replaced by ADD_11602

//ADD_7805 replaced by ADD_11601

//ADD_7804 replaced by ADD_11602

//ADD_7803 replaced by ADD_11602

//ADD_7802 replaced by ADD_11602

//ADD_7801 replaced by ADD_11602

//ADD_7809 replaced by ADD_11602

//ADD_7808 replaced by ADD_11602

//ADD_7807 replaced by ADD_11602

//ADD_7806 replaced by ADD_11602

//BADD_2593 replaced by BADD_2824

//BADD_2592 replaced by BADD_2823

//BADD_2591 replaced by BADD_2822

//ADD_7811 replaced by ADD_11602

//ADD_7810 replaced by ADD_11602

//KaratsubaCore_1244 replaced by KaratsubaCore_1437

//KaratsubaCore_1243 replaced by KaratsubaCore_1438

//KaratsubaCore_1242 replaced by KaratsubaCore_1437

//BADD_2597 replaced by BADD_2818

//BADD_2596 replaced by BADD_2820

//BADD_2595 replaced by BADD_2819

//BADD_2594 replaced by BADD_2818

//ADD_7813 replaced by ADD_8288

//ADD_7812 replaced by ADD_8288

//KaratsubaCore_1247 replaced by KaratsubaCore_1438

//KaratsubaCore_1246 replaced by KaratsubaCore_1435

//KaratsubaCore_1245 replaced by KaratsubaCore_1438

//BADD_2600 replaced by BADD_2824

//BADD_2599 replaced by BADD_2823

//BADD_2598 replaced by BADD_2822

//ADD_7815 replaced by ADD_11602

//ADD_7814 replaced by ADD_11602

//KaratsubaCore_1250 replaced by KaratsubaCore_1437

//KaratsubaCore_1249 replaced by KaratsubaCore_1438

//KaratsubaCore_1248 replaced by KaratsubaCore_1437

//ADD_7821 replaced by ADD_11602

//ADD_7820 replaced by ADD_11602

//ADD_7819 replaced by ADD_11602

//ADD_7818 replaced by ADD_11602

//ADD_7817 replaced by ADD_11602

//ADD_7816 replaced by ADD_11602

//ADD_7826 replaced by ADD_11601

//ADD_7825 replaced by ADD_11602

//ADD_7824 replaced by ADD_11602

//ADD_7823 replaced by ADD_11602

//ADD_7822 replaced by ADD_11602

//ADD_7830 replaced by ADD_11602

//ADD_7829 replaced by ADD_11602

//ADD_7828 replaced by ADD_11602

//ADD_7827 replaced by ADD_11602

//BADD_2603 replaced by BADD_2824

//BADD_2602 replaced by BADD_2823

//BADD_2601 replaced by BADD_2822

//ADD_7832 replaced by ADD_11602

//ADD_7831 replaced by ADD_11602

//KaratsubaCore_1253 replaced by KaratsubaCore_1437

//KaratsubaCore_1252 replaced by KaratsubaCore_1438

//KaratsubaCore_1251 replaced by KaratsubaCore_1437

//BADD_2607 replaced by BADD_2818

//BADD_2606 replaced by BADD_2820

//BADD_2605 replaced by BADD_2819

//BADD_2604 replaced by BADD_2818

//ADD_7834 replaced by ADD_8288

//ADD_7833 replaced by ADD_8288

//KaratsubaCore_1256 replaced by KaratsubaCore_1438

//KaratsubaCore_1255 replaced by KaratsubaCore_1435

//KaratsubaCore_1254 replaced by KaratsubaCore_1438

//BADD_2610 replaced by BADD_2824

//BADD_2609 replaced by BADD_2823

//BADD_2608 replaced by BADD_2822

//ADD_7836 replaced by ADD_11602

//ADD_7835 replaced by ADD_11602

//KaratsubaCore_1259 replaced by KaratsubaCore_1437

//KaratsubaCore_1258 replaced by KaratsubaCore_1438

//KaratsubaCore_1257 replaced by KaratsubaCore_1437

//ADD_7841 replaced by ADD_11595

//ADD_7840 replaced by ADD_11602

//ADD_7839 replaced by ADD_11602

//ADD_7838 replaced by ADD_11602

//ADD_7837 replaced by ADD_11602

//ADD_7846 replaced by ADD_11592

//ADD_7845 replaced by ADD_11602

//ADD_7844 replaced by ADD_11602

//ADD_7843 replaced by ADD_11602

//ADD_7842 replaced by ADD_11602

//ADD_7851 replaced by ADD_11592

//ADD_7850 replaced by ADD_11602

//ADD_7849 replaced by ADD_11602

//ADD_7848 replaced by ADD_11602

//ADD_7847 replaced by ADD_11602

//ADD_7856 replaced by ADD_11595

//ADD_7855 replaced by ADD_11602

//ADD_7854 replaced by ADD_11602

//ADD_7853 replaced by ADD_11602

//ADD_7852 replaced by ADD_11602

//BADD_2614 replaced by BADD_2818

//BADD_2613 replaced by BADD_2820

//BADD_2612 replaced by BADD_2819

//BADD_2611 replaced by BADD_2818

//ADD_7858 replaced by ADD_8288

//ADD_7857 replaced by ADD_8288

//KaratsubaCore_1262 replaced by KaratsubaCore_1438

//KaratsubaCore_1261 replaced by KaratsubaCore_1435

//KaratsubaCore_1260 replaced by KaratsubaCore_1438

//BADD_2618 replaced by BADD_2807

//BADD_2617 replaced by BADD_2809

//BADD_2616 replaced by BADD_2808

//BADD_2615 replaced by BADD_2807

//ADD_7860 replaced by ADD_8267

//ADD_7859 replaced by ADD_8267

//KaratsubaCore_1265 replaced by KaratsubaCore_1435

//KaratsubaCore_1264 replaced by KaratsubaCore_1426

//KaratsubaCore_1263 replaced by KaratsubaCore_1435

//BADD_2622 replaced by BADD_2818

//BADD_2621 replaced by BADD_2820

//BADD_2620 replaced by BADD_2819

//BADD_2619 replaced by BADD_2818

//ADD_7862 replaced by ADD_8288

//ADD_7861 replaced by ADD_8288

//KaratsubaCore_1268 replaced by KaratsubaCore_1438

//KaratsubaCore_1267 replaced by KaratsubaCore_1435

//KaratsubaCore_1266 replaced by KaratsubaCore_1438

//ADD_7868 replaced by ADD_11602

//ADD_7867 replaced by ADD_11602

//ADD_7866 replaced by ADD_11602

//ADD_7865 replaced by ADD_11602

//ADD_7864 replaced by ADD_11602

//ADD_7863 replaced by ADD_11602

//ADD_7873 replaced by ADD_11601

//ADD_7872 replaced by ADD_11602

//ADD_7871 replaced by ADD_11602

//ADD_7870 replaced by ADD_11602

//ADD_7869 replaced by ADD_11602

//ADD_7877 replaced by ADD_11602

//ADD_7876 replaced by ADD_11602

//ADD_7875 replaced by ADD_11602

//ADD_7874 replaced by ADD_11602

//BADD_2625 replaced by BADD_2824

//BADD_2624 replaced by BADD_2823

//BADD_2623 replaced by BADD_2822

//ADD_7879 replaced by ADD_11602

//ADD_7878 replaced by ADD_11602

//KaratsubaCore_1271 replaced by KaratsubaCore_1437

//KaratsubaCore_1270 replaced by KaratsubaCore_1438

//KaratsubaCore_1269 replaced by KaratsubaCore_1437

//BADD_2629 replaced by BADD_2818

//BADD_2628 replaced by BADD_2820

//BADD_2627 replaced by BADD_2819

//BADD_2626 replaced by BADD_2818

//ADD_7881 replaced by ADD_8288

//ADD_7880 replaced by ADD_8288

//KaratsubaCore_1274 replaced by KaratsubaCore_1438

//KaratsubaCore_1273 replaced by KaratsubaCore_1435

//KaratsubaCore_1272 replaced by KaratsubaCore_1438

//BADD_2632 replaced by BADD_2824

//BADD_2631 replaced by BADD_2823

//BADD_2630 replaced by BADD_2822

//ADD_7883 replaced by ADD_11602

//ADD_7882 replaced by ADD_11602

//KaratsubaCore_1277 replaced by KaratsubaCore_1437

//KaratsubaCore_1276 replaced by KaratsubaCore_1438

//KaratsubaCore_1275 replaced by KaratsubaCore_1437

//ADD_7889 replaced by ADD_11602

//ADD_7888 replaced by ADD_11602

//ADD_7887 replaced by ADD_11602

//ADD_7886 replaced by ADD_11602

//ADD_7885 replaced by ADD_11602

//ADD_7884 replaced by ADD_11602

//ADD_7894 replaced by ADD_11601

//ADD_7893 replaced by ADD_11602

//ADD_7892 replaced by ADD_11602

//ADD_7891 replaced by ADD_11602

//ADD_7890 replaced by ADD_11602

//ADD_7898 replaced by ADD_11602

//ADD_7897 replaced by ADD_11602

//ADD_7896 replaced by ADD_11602

//ADD_7895 replaced by ADD_11602

//BADD_2635 replaced by BADD_2824

//BADD_2634 replaced by BADD_2823

//BADD_2633 replaced by BADD_2822

//ADD_7900 replaced by ADD_11602

//ADD_7899 replaced by ADD_11602

//KaratsubaCore_1280 replaced by KaratsubaCore_1437

//KaratsubaCore_1279 replaced by KaratsubaCore_1438

//KaratsubaCore_1278 replaced by KaratsubaCore_1437

//BADD_2639 replaced by BADD_2818

//BADD_2638 replaced by BADD_2820

//BADD_2637 replaced by BADD_2819

//BADD_2636 replaced by BADD_2818

//ADD_7902 replaced by ADD_8288

//ADD_7901 replaced by ADD_8288

//KaratsubaCore_1283 replaced by KaratsubaCore_1438

//KaratsubaCore_1282 replaced by KaratsubaCore_1435

//KaratsubaCore_1281 replaced by KaratsubaCore_1438

//BADD_2642 replaced by BADD_2824

//BADD_2641 replaced by BADD_2823

//BADD_2640 replaced by BADD_2822

//ADD_7904 replaced by ADD_11602

//ADD_7903 replaced by ADD_11602

//KaratsubaCore_1286 replaced by KaratsubaCore_1437

//KaratsubaCore_1285 replaced by KaratsubaCore_1438

//KaratsubaCore_1284 replaced by KaratsubaCore_1437

//ADD_7909 replaced by ADD_11595

//ADD_7908 replaced by ADD_11602

//ADD_7907 replaced by ADD_11602

//ADD_7906 replaced by ADD_11602

//ADD_7905 replaced by ADD_11602

//ADD_7914 replaced by ADD_11592

//ADD_7913 replaced by ADD_11602

//ADD_7912 replaced by ADD_11602

//ADD_7911 replaced by ADD_11602

//ADD_7910 replaced by ADD_11602

//ADD_7919 replaced by ADD_11592

//ADD_7918 replaced by ADD_11602

//ADD_7917 replaced by ADD_11602

//ADD_7916 replaced by ADD_11602

//ADD_7915 replaced by ADD_11602

//ADD_7924 replaced by ADD_11595

//ADD_7923 replaced by ADD_11602

//ADD_7922 replaced by ADD_11602

//ADD_7921 replaced by ADD_11602

//ADD_7920 replaced by ADD_11602

//BADD_2646 replaced by BADD_2818

//BADD_2645 replaced by BADD_2820

//BADD_2644 replaced by BADD_2819

//BADD_2643 replaced by BADD_2818

//ADD_7926 replaced by ADD_8288

//ADD_7925 replaced by ADD_8288

//KaratsubaCore_1289 replaced by KaratsubaCore_1438

//KaratsubaCore_1288 replaced by KaratsubaCore_1435

//KaratsubaCore_1287 replaced by KaratsubaCore_1438

//BADD_2650 replaced by BADD_2807

//BADD_2649 replaced by BADD_2809

//BADD_2648 replaced by BADD_2808

//BADD_2647 replaced by BADD_2807

//ADD_7928 replaced by ADD_8267

//ADD_7927 replaced by ADD_8267

//KaratsubaCore_1292 replaced by KaratsubaCore_1435

//KaratsubaCore_1291 replaced by KaratsubaCore_1426

//KaratsubaCore_1290 replaced by KaratsubaCore_1435

//BADD_2654 replaced by BADD_2818

//BADD_2653 replaced by BADD_2820

//BADD_2652 replaced by BADD_2819

//BADD_2651 replaced by BADD_2818

//ADD_7930 replaced by ADD_8288

//ADD_7929 replaced by ADD_8288

//KaratsubaCore_1295 replaced by KaratsubaCore_1438

//KaratsubaCore_1294 replaced by KaratsubaCore_1435

//KaratsubaCore_1293 replaced by KaratsubaCore_1438

//ADD_7936 replaced by ADD_11602

//ADD_7935 replaced by ADD_11602

//ADD_7934 replaced by ADD_11602

//ADD_7933 replaced by ADD_11602

//ADD_7932 replaced by ADD_11602

//ADD_7931 replaced by ADD_11602

//ADD_7941 replaced by ADD_11601

//ADD_7940 replaced by ADD_11602

//ADD_7939 replaced by ADD_11602

//ADD_7938 replaced by ADD_11602

//ADD_7937 replaced by ADD_11602

//ADD_7945 replaced by ADD_11602

//ADD_7944 replaced by ADD_11602

//ADD_7943 replaced by ADD_11602

//ADD_7942 replaced by ADD_11602

//BADD_2657 replaced by BADD_2824

//BADD_2656 replaced by BADD_2823

//BADD_2655 replaced by BADD_2822

//ADD_7947 replaced by ADD_11602

//ADD_7946 replaced by ADD_11602

//KaratsubaCore_1298 replaced by KaratsubaCore_1437

//KaratsubaCore_1297 replaced by KaratsubaCore_1438

//KaratsubaCore_1296 replaced by KaratsubaCore_1437

//BADD_2661 replaced by BADD_2818

//BADD_2660 replaced by BADD_2820

//BADD_2659 replaced by BADD_2819

//BADD_2658 replaced by BADD_2818

//ADD_7949 replaced by ADD_8288

//ADD_7948 replaced by ADD_8288

//KaratsubaCore_1301 replaced by KaratsubaCore_1438

//KaratsubaCore_1300 replaced by KaratsubaCore_1435

//KaratsubaCore_1299 replaced by KaratsubaCore_1438

//BADD_2664 replaced by BADD_2824

//BADD_2663 replaced by BADD_2823

//BADD_2662 replaced by BADD_2822

//ADD_7951 replaced by ADD_11602

//ADD_7950 replaced by ADD_11602

//KaratsubaCore_1304 replaced by KaratsubaCore_1437

//KaratsubaCore_1303 replaced by KaratsubaCore_1438

//KaratsubaCore_1302 replaced by KaratsubaCore_1437

//ADD_7957 replaced by ADD_11602

//ADD_7956 replaced by ADD_11602

//ADD_7955 replaced by ADD_11602

//ADD_7954 replaced by ADD_11602

//ADD_7953 replaced by ADD_11602

//ADD_7952 replaced by ADD_11602

//ADD_7962 replaced by ADD_11601

//ADD_7961 replaced by ADD_11602

//ADD_7960 replaced by ADD_11602

//ADD_7959 replaced by ADD_11602

//ADD_7958 replaced by ADD_11602

//ADD_7966 replaced by ADD_11602

//ADD_7965 replaced by ADD_11602

//ADD_7964 replaced by ADD_11602

//ADD_7963 replaced by ADD_11602

//BADD_2667 replaced by BADD_2824

//BADD_2666 replaced by BADD_2823

//BADD_2665 replaced by BADD_2822

//ADD_7968 replaced by ADD_11602

//ADD_7967 replaced by ADD_11602

//KaratsubaCore_1307 replaced by KaratsubaCore_1437

//KaratsubaCore_1306 replaced by KaratsubaCore_1438

//KaratsubaCore_1305 replaced by KaratsubaCore_1437

//BADD_2671 replaced by BADD_2818

//BADD_2670 replaced by BADD_2820

//BADD_2669 replaced by BADD_2819

//BADD_2668 replaced by BADD_2818

//ADD_7970 replaced by ADD_8288

//ADD_7969 replaced by ADD_8288

//KaratsubaCore_1310 replaced by KaratsubaCore_1438

//KaratsubaCore_1309 replaced by KaratsubaCore_1435

//KaratsubaCore_1308 replaced by KaratsubaCore_1438

//BADD_2674 replaced by BADD_2824

//BADD_2673 replaced by BADD_2823

//BADD_2672 replaced by BADD_2822

//ADD_7972 replaced by ADD_11602

//ADD_7971 replaced by ADD_11602

//KaratsubaCore_1313 replaced by KaratsubaCore_1437

//KaratsubaCore_1312 replaced by KaratsubaCore_1438

//KaratsubaCore_1311 replaced by KaratsubaCore_1437

//ADD_7977 replaced by ADD_11595

//ADD_7976 replaced by ADD_11602

//ADD_7975 replaced by ADD_11602

//ADD_7974 replaced by ADD_11602

//ADD_7973 replaced by ADD_11602

//ADD_7982 replaced by ADD_11592

//ADD_7981 replaced by ADD_11602

//ADD_7980 replaced by ADD_11602

//ADD_7979 replaced by ADD_11602

//ADD_7978 replaced by ADD_11602

//ADD_7987 replaced by ADD_11592

//ADD_7986 replaced by ADD_11602

//ADD_7985 replaced by ADD_11602

//ADD_7984 replaced by ADD_11602

//ADD_7983 replaced by ADD_11602

//ADD_7992 replaced by ADD_11595

//ADD_7991 replaced by ADD_11602

//ADD_7990 replaced by ADD_11602

//ADD_7989 replaced by ADD_11602

//ADD_7988 replaced by ADD_11602

//BADD_2678 replaced by BADD_2818

//BADD_2677 replaced by BADD_2820

//BADD_2676 replaced by BADD_2819

//BADD_2675 replaced by BADD_2818

//ADD_7994 replaced by ADD_8288

//ADD_7993 replaced by ADD_8288

//KaratsubaCore_1316 replaced by KaratsubaCore_1438

//KaratsubaCore_1315 replaced by KaratsubaCore_1435

//KaratsubaCore_1314 replaced by KaratsubaCore_1438

//BADD_2682 replaced by BADD_2807

//BADD_2681 replaced by BADD_2809

//BADD_2680 replaced by BADD_2808

//BADD_2679 replaced by BADD_2807

//ADD_7996 replaced by ADD_8267

//ADD_7995 replaced by ADD_8267

//KaratsubaCore_1319 replaced by KaratsubaCore_1435

//KaratsubaCore_1318 replaced by KaratsubaCore_1426

//KaratsubaCore_1317 replaced by KaratsubaCore_1435

//BADD_2686 replaced by BADD_2818

//BADD_2685 replaced by BADD_2820

//BADD_2684 replaced by BADD_2819

//BADD_2683 replaced by BADD_2818

//ADD_7998 replaced by ADD_8288

//ADD_7997 replaced by ADD_8288

//KaratsubaCore_1322 replaced by KaratsubaCore_1438

//KaratsubaCore_1321 replaced by KaratsubaCore_1435

//KaratsubaCore_1320 replaced by KaratsubaCore_1438

//ADD_8004 replaced by ADD_11602

//ADD_8003 replaced by ADD_11602

//ADD_8002 replaced by ADD_11602

//ADD_8001 replaced by ADD_11602

//ADD_8000 replaced by ADD_11602

//ADD_7999 replaced by ADD_11602

//ADD_8009 replaced by ADD_11601

//ADD_8008 replaced by ADD_11602

//ADD_8007 replaced by ADD_11602

//ADD_8006 replaced by ADD_11602

//ADD_8005 replaced by ADD_11602

//ADD_8013 replaced by ADD_11602

//ADD_8012 replaced by ADD_11602

//ADD_8011 replaced by ADD_11602

//ADD_8010 replaced by ADD_11602

//BADD_2689 replaced by BADD_2824

//BADD_2688 replaced by BADD_2823

//BADD_2687 replaced by BADD_2822

//ADD_8015 replaced by ADD_11602

//ADD_8014 replaced by ADD_11602

//KaratsubaCore_1325 replaced by KaratsubaCore_1437

//KaratsubaCore_1324 replaced by KaratsubaCore_1438

//KaratsubaCore_1323 replaced by KaratsubaCore_1437

//BADD_2693 replaced by BADD_2818

//BADD_2692 replaced by BADD_2820

//BADD_2691 replaced by BADD_2819

//BADD_2690 replaced by BADD_2818

//ADD_8017 replaced by ADD_8288

//ADD_8016 replaced by ADD_8288

//KaratsubaCore_1328 replaced by KaratsubaCore_1438

//KaratsubaCore_1327 replaced by KaratsubaCore_1435

//KaratsubaCore_1326 replaced by KaratsubaCore_1438

//BADD_2696 replaced by BADD_2824

//BADD_2695 replaced by BADD_2823

//BADD_2694 replaced by BADD_2822

//ADD_8019 replaced by ADD_11602

//ADD_8018 replaced by ADD_11602

//KaratsubaCore_1331 replaced by KaratsubaCore_1437

//KaratsubaCore_1330 replaced by KaratsubaCore_1438

//KaratsubaCore_1329 replaced by KaratsubaCore_1437

//ADD_8025 replaced by ADD_11602

//ADD_8024 replaced by ADD_11602

//ADD_8023 replaced by ADD_11602

//ADD_8022 replaced by ADD_11602

//ADD_8021 replaced by ADD_11602

//ADD_8020 replaced by ADD_11602

//ADD_8030 replaced by ADD_11601

//ADD_8029 replaced by ADD_11602

//ADD_8028 replaced by ADD_11602

//ADD_8027 replaced by ADD_11602

//ADD_8026 replaced by ADD_11602

//ADD_8034 replaced by ADD_11602

//ADD_8033 replaced by ADD_11602

//ADD_8032 replaced by ADD_11602

//ADD_8031 replaced by ADD_11602

//BADD_2699 replaced by BADD_2824

//BADD_2698 replaced by BADD_2823

//BADD_2697 replaced by BADD_2822

//ADD_8036 replaced by ADD_11602

//ADD_8035 replaced by ADD_11602

//KaratsubaCore_1334 replaced by KaratsubaCore_1437

//KaratsubaCore_1333 replaced by KaratsubaCore_1438

//KaratsubaCore_1332 replaced by KaratsubaCore_1437

//BADD_2703 replaced by BADD_2818

//BADD_2702 replaced by BADD_2820

//BADD_2701 replaced by BADD_2819

//BADD_2700 replaced by BADD_2818

//ADD_8038 replaced by ADD_8288

//ADD_8037 replaced by ADD_8288

//KaratsubaCore_1337 replaced by KaratsubaCore_1438

//KaratsubaCore_1336 replaced by KaratsubaCore_1435

//KaratsubaCore_1335 replaced by KaratsubaCore_1438

//BADD_2706 replaced by BADD_2824

//BADD_2705 replaced by BADD_2823

//BADD_2704 replaced by BADD_2822

//ADD_8040 replaced by ADD_11602

//ADD_8039 replaced by ADD_11602

//KaratsubaCore_1340 replaced by KaratsubaCore_1437

//KaratsubaCore_1339 replaced by KaratsubaCore_1438

//KaratsubaCore_1338 replaced by KaratsubaCore_1437

//ADD_8045 replaced by ADD_11595

//ADD_8044 replaced by ADD_11602

//ADD_8043 replaced by ADD_11602

//ADD_8042 replaced by ADD_11602

//ADD_8041 replaced by ADD_11602

//ADD_8050 replaced by ADD_11592

//ADD_8049 replaced by ADD_11602

//ADD_8048 replaced by ADD_11602

//ADD_8047 replaced by ADD_11602

//ADD_8046 replaced by ADD_11602

//ADD_8055 replaced by ADD_11592

//ADD_8054 replaced by ADD_11602

//ADD_8053 replaced by ADD_11602

//ADD_8052 replaced by ADD_11602

//ADD_8051 replaced by ADD_11602

//ADD_8060 replaced by ADD_11595

//ADD_8059 replaced by ADD_11602

//ADD_8058 replaced by ADD_11602

//ADD_8057 replaced by ADD_11602

//ADD_8056 replaced by ADD_11602

//BADD_2710 replaced by BADD_2818

//BADD_2709 replaced by BADD_2820

//BADD_2708 replaced by BADD_2819

//BADD_2707 replaced by BADD_2818

//ADD_8062 replaced by ADD_8288

//ADD_8061 replaced by ADD_8288

//KaratsubaCore_1343 replaced by KaratsubaCore_1438

//KaratsubaCore_1342 replaced by KaratsubaCore_1435

//KaratsubaCore_1341 replaced by KaratsubaCore_1438

//BADD_2714 replaced by BADD_2807

//BADD_2713 replaced by BADD_2809

//BADD_2712 replaced by BADD_2808

//BADD_2711 replaced by BADD_2807

//ADD_8064 replaced by ADD_8267

//ADD_8063 replaced by ADD_8267

//KaratsubaCore_1346 replaced by KaratsubaCore_1435

//KaratsubaCore_1345 replaced by KaratsubaCore_1426

//KaratsubaCore_1344 replaced by KaratsubaCore_1435

//BADD_2718 replaced by BADD_2818

//BADD_2717 replaced by BADD_2820

//BADD_2716 replaced by BADD_2819

//BADD_2715 replaced by BADD_2818

//ADD_8066 replaced by ADD_8288

//ADD_8065 replaced by ADD_8288

//KaratsubaCore_1349 replaced by KaratsubaCore_1438

//KaratsubaCore_1348 replaced by KaratsubaCore_1435

//KaratsubaCore_1347 replaced by KaratsubaCore_1438

//ADD_8072 replaced by ADD_11602

//ADD_8071 replaced by ADD_11602

//ADD_8070 replaced by ADD_11602

//ADD_8069 replaced by ADD_11602

//ADD_8068 replaced by ADD_11602

//ADD_8067 replaced by ADD_11602

//ADD_8077 replaced by ADD_11601

//ADD_8076 replaced by ADD_11602

//ADD_8075 replaced by ADD_11602

//ADD_8074 replaced by ADD_11602

//ADD_8073 replaced by ADD_11602

//ADD_8081 replaced by ADD_11602

//ADD_8080 replaced by ADD_11602

//ADD_8079 replaced by ADD_11602

//ADD_8078 replaced by ADD_11602

//BADD_2721 replaced by BADD_2824

//BADD_2720 replaced by BADD_2823

//BADD_2719 replaced by BADD_2822

//ADD_8083 replaced by ADD_11602

//ADD_8082 replaced by ADD_11602

//KaratsubaCore_1352 replaced by KaratsubaCore_1437

//KaratsubaCore_1351 replaced by KaratsubaCore_1438

//KaratsubaCore_1350 replaced by KaratsubaCore_1437

//BADD_2725 replaced by BADD_2818

//BADD_2724 replaced by BADD_2820

//BADD_2723 replaced by BADD_2819

//BADD_2722 replaced by BADD_2818

//ADD_8085 replaced by ADD_8288

//ADD_8084 replaced by ADD_8288

//KaratsubaCore_1355 replaced by KaratsubaCore_1438

//KaratsubaCore_1354 replaced by KaratsubaCore_1435

//KaratsubaCore_1353 replaced by KaratsubaCore_1438

//BADD_2728 replaced by BADD_2824

//BADD_2727 replaced by BADD_2823

//BADD_2726 replaced by BADD_2822

//ADD_8087 replaced by ADD_11602

//ADD_8086 replaced by ADD_11602

//KaratsubaCore_1358 replaced by KaratsubaCore_1437

//KaratsubaCore_1357 replaced by KaratsubaCore_1438

//KaratsubaCore_1356 replaced by KaratsubaCore_1437

//ADD_8093 replaced by ADD_11602

//ADD_8092 replaced by ADD_11602

//ADD_8091 replaced by ADD_11602

//ADD_8090 replaced by ADD_11602

//ADD_8089 replaced by ADD_11602

//ADD_8088 replaced by ADD_11602

//ADD_8098 replaced by ADD_11601

//ADD_8097 replaced by ADD_11602

//ADD_8096 replaced by ADD_11602

//ADD_8095 replaced by ADD_11602

//ADD_8094 replaced by ADD_11602

//ADD_8102 replaced by ADD_11602

//ADD_8101 replaced by ADD_11602

//ADD_8100 replaced by ADD_11602

//ADD_8099 replaced by ADD_11602

//BADD_2731 replaced by BADD_2824

//BADD_2730 replaced by BADD_2823

//BADD_2729 replaced by BADD_2822

//ADD_8104 replaced by ADD_11602

//ADD_8103 replaced by ADD_11602

//KaratsubaCore_1361 replaced by KaratsubaCore_1437

//KaratsubaCore_1360 replaced by KaratsubaCore_1438

//KaratsubaCore_1359 replaced by KaratsubaCore_1437

//BADD_2735 replaced by BADD_2818

//BADD_2734 replaced by BADD_2820

//BADD_2733 replaced by BADD_2819

//BADD_2732 replaced by BADD_2818

//ADD_8106 replaced by ADD_8288

//ADD_8105 replaced by ADD_8288

//KaratsubaCore_1364 replaced by KaratsubaCore_1438

//KaratsubaCore_1363 replaced by KaratsubaCore_1435

//KaratsubaCore_1362 replaced by KaratsubaCore_1438

//BADD_2738 replaced by BADD_2824

//BADD_2737 replaced by BADD_2823

//BADD_2736 replaced by BADD_2822

//ADD_8108 replaced by ADD_11602

//ADD_8107 replaced by ADD_11602

//KaratsubaCore_1367 replaced by KaratsubaCore_1437

//KaratsubaCore_1366 replaced by KaratsubaCore_1438

//KaratsubaCore_1365 replaced by KaratsubaCore_1437

//ADD_8113 replaced by ADD_11595

//ADD_8112 replaced by ADD_11602

//ADD_8111 replaced by ADD_11602

//ADD_8110 replaced by ADD_11602

//ADD_8109 replaced by ADD_11602

//ADD_8118 replaced by ADD_11592

//ADD_8117 replaced by ADD_11602

//ADD_8116 replaced by ADD_11602

//ADD_8115 replaced by ADD_11602

//ADD_8114 replaced by ADD_11602

//ADD_8123 replaced by ADD_11592

//ADD_8122 replaced by ADD_11602

//ADD_8121 replaced by ADD_11602

//ADD_8120 replaced by ADD_11602

//ADD_8119 replaced by ADD_11602

//ADD_8128 replaced by ADD_11595

//ADD_8127 replaced by ADD_11602

//ADD_8126 replaced by ADD_11602

//ADD_8125 replaced by ADD_11602

//ADD_8124 replaced by ADD_11602

//BADD_2742 replaced by BADD_2818

//BADD_2741 replaced by BADD_2820

//BADD_2740 replaced by BADD_2819

//BADD_2739 replaced by BADD_2818

//ADD_8130 replaced by ADD_8288

//ADD_8129 replaced by ADD_8288

//KaratsubaCore_1370 replaced by KaratsubaCore_1438

//KaratsubaCore_1369 replaced by KaratsubaCore_1435

//KaratsubaCore_1368 replaced by KaratsubaCore_1438

//BADD_2746 replaced by BADD_2807

//BADD_2745 replaced by BADD_2809

//BADD_2744 replaced by BADD_2808

//BADD_2743 replaced by BADD_2807

//ADD_8132 replaced by ADD_8267

//ADD_8131 replaced by ADD_8267

//KaratsubaCore_1373 replaced by KaratsubaCore_1435

//KaratsubaCore_1372 replaced by KaratsubaCore_1426

//KaratsubaCore_1371 replaced by KaratsubaCore_1435

//BADD_2750 replaced by BADD_2818

//BADD_2749 replaced by BADD_2820

//BADD_2748 replaced by BADD_2819

//BADD_2747 replaced by BADD_2818

//ADD_8134 replaced by ADD_8288

//ADD_8133 replaced by ADD_8288

//KaratsubaCore_1376 replaced by KaratsubaCore_1438

//KaratsubaCore_1375 replaced by KaratsubaCore_1435

//KaratsubaCore_1374 replaced by KaratsubaCore_1438

//ADD_8140 replaced by ADD_11602

//ADD_8139 replaced by ADD_11602

//ADD_8138 replaced by ADD_11602

//ADD_8137 replaced by ADD_11602

//ADD_8136 replaced by ADD_11602

//ADD_8135 replaced by ADD_11602

//ADD_8145 replaced by ADD_11601

//ADD_8144 replaced by ADD_11602

//ADD_8143 replaced by ADD_11602

//ADD_8142 replaced by ADD_11602

//ADD_8141 replaced by ADD_11602

//ADD_8149 replaced by ADD_11602

//ADD_8148 replaced by ADD_11602

//ADD_8147 replaced by ADD_11602

//ADD_8146 replaced by ADD_11602

//BADD_2753 replaced by BADD_2824

//BADD_2752 replaced by BADD_2823

//BADD_2751 replaced by BADD_2822

//ADD_8151 replaced by ADD_11602

//ADD_8150 replaced by ADD_11602

//KaratsubaCore_1379 replaced by KaratsubaCore_1437

//KaratsubaCore_1378 replaced by KaratsubaCore_1438

//KaratsubaCore_1377 replaced by KaratsubaCore_1437

//BADD_2757 replaced by BADD_2818

//BADD_2756 replaced by BADD_2820

//BADD_2755 replaced by BADD_2819

//BADD_2754 replaced by BADD_2818

//ADD_8153 replaced by ADD_8288

//ADD_8152 replaced by ADD_8288

//KaratsubaCore_1382 replaced by KaratsubaCore_1438

//KaratsubaCore_1381 replaced by KaratsubaCore_1435

//KaratsubaCore_1380 replaced by KaratsubaCore_1438

//BADD_2760 replaced by BADD_2824

//BADD_2759 replaced by BADD_2823

//BADD_2758 replaced by BADD_2822

//ADD_8155 replaced by ADD_11602

//ADD_8154 replaced by ADD_11602

//KaratsubaCore_1385 replaced by KaratsubaCore_1437

//KaratsubaCore_1384 replaced by KaratsubaCore_1438

//KaratsubaCore_1383 replaced by KaratsubaCore_1437

//ADD_8161 replaced by ADD_11602

//ADD_8160 replaced by ADD_11602

//ADD_8159 replaced by ADD_11602

//ADD_8158 replaced by ADD_11602

//ADD_8157 replaced by ADD_11602

//ADD_8156 replaced by ADD_11602

//ADD_8166 replaced by ADD_11601

//ADD_8165 replaced by ADD_11602

//ADD_8164 replaced by ADD_11602

//ADD_8163 replaced by ADD_11602

//ADD_8162 replaced by ADD_11602

//ADD_8170 replaced by ADD_11602

//ADD_8169 replaced by ADD_11602

//ADD_8168 replaced by ADD_11602

//ADD_8167 replaced by ADD_11602

//BADD_2763 replaced by BADD_2824

//BADD_2762 replaced by BADD_2823

//BADD_2761 replaced by BADD_2822

//ADD_8172 replaced by ADD_11602

//ADD_8171 replaced by ADD_11602

//KaratsubaCore_1388 replaced by KaratsubaCore_1437

//KaratsubaCore_1387 replaced by KaratsubaCore_1438

//KaratsubaCore_1386 replaced by KaratsubaCore_1437

//BADD_2767 replaced by BADD_2818

//BADD_2766 replaced by BADD_2820

//BADD_2765 replaced by BADD_2819

//BADD_2764 replaced by BADD_2818

//ADD_8174 replaced by ADD_8288

//ADD_8173 replaced by ADD_8288

//KaratsubaCore_1391 replaced by KaratsubaCore_1438

//KaratsubaCore_1390 replaced by KaratsubaCore_1435

//KaratsubaCore_1389 replaced by KaratsubaCore_1438

//BADD_2770 replaced by BADD_2824

//BADD_2769 replaced by BADD_2823

//BADD_2768 replaced by BADD_2822

//ADD_8176 replaced by ADD_11602

//ADD_8175 replaced by ADD_11602

//KaratsubaCore_1394 replaced by KaratsubaCore_1437

//KaratsubaCore_1393 replaced by KaratsubaCore_1438

//KaratsubaCore_1392 replaced by KaratsubaCore_1437

//ADD_8181 replaced by ADD_11595

//ADD_8180 replaced by ADD_11602

//ADD_8179 replaced by ADD_11602

//ADD_8178 replaced by ADD_11602

//ADD_8177 replaced by ADD_11602

//ADD_8186 replaced by ADD_11592

//ADD_8185 replaced by ADD_11602

//ADD_8184 replaced by ADD_11602

//ADD_8183 replaced by ADD_11602

//ADD_8182 replaced by ADD_11602

//ADD_8191 replaced by ADD_11592

//ADD_8190 replaced by ADD_11602

//ADD_8189 replaced by ADD_11602

//ADD_8188 replaced by ADD_11602

//ADD_8187 replaced by ADD_11602

//ADD_8196 replaced by ADD_11595

//ADD_8195 replaced by ADD_11602

//ADD_8194 replaced by ADD_11602

//ADD_8193 replaced by ADD_11602

//ADD_8192 replaced by ADD_11602

//BADD_2774 replaced by BADD_2818

//BADD_2773 replaced by BADD_2820

//BADD_2772 replaced by BADD_2819

//BADD_2771 replaced by BADD_2818

//ADD_8198 replaced by ADD_8288

//ADD_8197 replaced by ADD_8288

//KaratsubaCore_1397 replaced by KaratsubaCore_1438

//KaratsubaCore_1396 replaced by KaratsubaCore_1435

//KaratsubaCore_1395 replaced by KaratsubaCore_1438

//BADD_2778 replaced by BADD_2807

//BADD_2777 replaced by BADD_2809

//BADD_2776 replaced by BADD_2808

//BADD_2775 replaced by BADD_2807

//ADD_8200 replaced by ADD_8267

//ADD_8199 replaced by ADD_8267

//KaratsubaCore_1400 replaced by KaratsubaCore_1435

//KaratsubaCore_1399 replaced by KaratsubaCore_1426

//KaratsubaCore_1398 replaced by KaratsubaCore_1435

//BADD_2782 replaced by BADD_2818

//BADD_2781 replaced by BADD_2820

//BADD_2780 replaced by BADD_2819

//BADD_2779 replaced by BADD_2818

//ADD_8202 replaced by ADD_8288

//ADD_8201 replaced by ADD_8288

//KaratsubaCore_1403 replaced by KaratsubaCore_1438

//KaratsubaCore_1402 replaced by KaratsubaCore_1435

//KaratsubaCore_1401 replaced by KaratsubaCore_1438

//ADD_8208 replaced by ADD_11602

//ADD_8207 replaced by ADD_11602

//ADD_8206 replaced by ADD_11602

//ADD_8205 replaced by ADD_11602

//ADD_8204 replaced by ADD_11602

//ADD_8203 replaced by ADD_11602

//ADD_8213 replaced by ADD_11601

//ADD_8212 replaced by ADD_11602

//ADD_8211 replaced by ADD_11602

//ADD_8210 replaced by ADD_11602

//ADD_8209 replaced by ADD_11602

//ADD_8217 replaced by ADD_11602

//ADD_8216 replaced by ADD_11602

//ADD_8215 replaced by ADD_11602

//ADD_8214 replaced by ADD_11602

//BADD_2785 replaced by BADD_2824

//BADD_2784 replaced by BADD_2823

//BADD_2783 replaced by BADD_2822

//ADD_8219 replaced by ADD_11602

//ADD_8218 replaced by ADD_11602

//KaratsubaCore_1406 replaced by KaratsubaCore_1437

//KaratsubaCore_1405 replaced by KaratsubaCore_1438

//KaratsubaCore_1404 replaced by KaratsubaCore_1437

//BADD_2789 replaced by BADD_2818

//BADD_2788 replaced by BADD_2820

//BADD_2787 replaced by BADD_2819

//BADD_2786 replaced by BADD_2818

//ADD_8221 replaced by ADD_8288

//ADD_8220 replaced by ADD_8288

//KaratsubaCore_1409 replaced by KaratsubaCore_1438

//KaratsubaCore_1408 replaced by KaratsubaCore_1435

//KaratsubaCore_1407 replaced by KaratsubaCore_1438

//BADD_2792 replaced by BADD_2824

//BADD_2791 replaced by BADD_2823

//BADD_2790 replaced by BADD_2822

//ADD_8223 replaced by ADD_11602

//ADD_8222 replaced by ADD_11602

//KaratsubaCore_1412 replaced by KaratsubaCore_1437

//KaratsubaCore_1411 replaced by KaratsubaCore_1438

//KaratsubaCore_1410 replaced by KaratsubaCore_1437

//ADD_8229 replaced by ADD_11602

//ADD_8228 replaced by ADD_11602

//ADD_8227 replaced by ADD_11602

//ADD_8226 replaced by ADD_11602

//ADD_8225 replaced by ADD_11602

//ADD_8224 replaced by ADD_11602

//ADD_8234 replaced by ADD_11601

//ADD_8233 replaced by ADD_11602

//ADD_8232 replaced by ADD_11602

//ADD_8231 replaced by ADD_11602

//ADD_8230 replaced by ADD_11602

//ADD_8238 replaced by ADD_11602

//ADD_8237 replaced by ADD_11602

//ADD_8236 replaced by ADD_11602

//ADD_8235 replaced by ADD_11602

//BADD_2795 replaced by BADD_2824

//BADD_2794 replaced by BADD_2823

//BADD_2793 replaced by BADD_2822

//ADD_8240 replaced by ADD_11602

//ADD_8239 replaced by ADD_11602

//KaratsubaCore_1415 replaced by KaratsubaCore_1437

//KaratsubaCore_1414 replaced by KaratsubaCore_1438

//KaratsubaCore_1413 replaced by KaratsubaCore_1437

//BADD_2799 replaced by BADD_2818

//BADD_2798 replaced by BADD_2820

//BADD_2797 replaced by BADD_2819

//BADD_2796 replaced by BADD_2818

//ADD_8242 replaced by ADD_8288

//ADD_8241 replaced by ADD_8288

//KaratsubaCore_1418 replaced by KaratsubaCore_1438

//KaratsubaCore_1417 replaced by KaratsubaCore_1435

//KaratsubaCore_1416 replaced by KaratsubaCore_1438

//BADD_2802 replaced by BADD_2824

//BADD_2801 replaced by BADD_2823

//BADD_2800 replaced by BADD_2822

//ADD_8244 replaced by ADD_11602

//ADD_8243 replaced by ADD_11602

//KaratsubaCore_1421 replaced by KaratsubaCore_1437

//KaratsubaCore_1420 replaced by KaratsubaCore_1438

//KaratsubaCore_1419 replaced by KaratsubaCore_1437

//ADD_8249 replaced by ADD_11595

//ADD_8248 replaced by ADD_11602

//ADD_8247 replaced by ADD_11602

//ADD_8246 replaced by ADD_11602

//ADD_8245 replaced by ADD_11602

//ADD_8254 replaced by ADD_11592

//ADD_8253 replaced by ADD_11602

//ADD_8252 replaced by ADD_11602

//ADD_8251 replaced by ADD_11602

//ADD_8250 replaced by ADD_11602

//ADD_8259 replaced by ADD_11592

//ADD_8258 replaced by ADD_11602

//ADD_8257 replaced by ADD_11602

//ADD_8256 replaced by ADD_11602

//ADD_8255 replaced by ADD_11602

//ADD_8264 replaced by ADD_11595

//ADD_8263 replaced by ADD_11602

//ADD_8262 replaced by ADD_11602

//ADD_8261 replaced by ADD_11602

//ADD_8260 replaced by ADD_11602

//BADD_2806 replaced by BADD_2818

//BADD_2805 replaced by BADD_2820

//BADD_2804 replaced by BADD_2819

//BADD_2803 replaced by BADD_2818

//ADD_8266 replaced by ADD_8288

//ADD_8265 replaced by ADD_8288

//KaratsubaCore_1424 replaced by KaratsubaCore_1438

//KaratsubaCore_1423 replaced by KaratsubaCore_1435

//KaratsubaCore_1422 replaced by KaratsubaCore_1438

//BADD_2810 replaced by BADD_2807

module BADD_2809 (
  input      [100:0]  io_a,
  input      [100:0]  io_b,
  input               io_c,
  output     [101:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [4:0]    adder_adds_2_io_A_0;
  wire       [4:0]    adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [5:0]    adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [4:0]    _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11560 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[4:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[4:0]), //i
    .io_CIN (_zz_io_CIN_1            ), //i
    .io_S   (adder_adds_2_io_S[5:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[100 : 96];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[100 : 96];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_s <= adder_adds_2_io_S[5];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[4 : 0];
  end


endmodule

module BADD_2808 (
  input      [100:0]  io_a,
  input      [100:0]  io_b,
  input               io_c,
  output     [101:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [4:0]    adder_adds_2_io_A_0;
  wire       [4:0]    adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [5:0]    adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [4:0]    _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11560 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[4:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[4:0]), //i
    .io_CIN (_zz_io_CIN_1            ), //i
    .io_S   (adder_adds_2_io_S[5:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[100 : 96];
  assign adder_adds_0_io_A_1 = (~ io_b[47 : 0]);
  assign adder_adds_1_io_A_1 = (~ io_b[95 : 48]);
  assign adder_adds_2_io_A_1 = (~ io_b[100 : 96]);
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_s <= (! adder_adds_2_io_S[5]);
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[4 : 0];
  end


endmodule

module BADD_2807 (
  input      [99:0]   io_a,
  input      [99:0]   io_b,
  input               io_c,
  output     [100:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [3:0]    adder_adds_2_io_A_0;
  wire       [3:0]    adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [4:0]    adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [3:0]    _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11563 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[3:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[3:0]), //i
    .io_CIN (_zz_io_CIN_1            ), //i
    .io_S   (adder_adds_2_io_S[4:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[99 : 96];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[99 : 96];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_s <= adder_adds_2_io_S[4];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[3 : 0];
  end


endmodule

//ADD_8268 replaced by ADD_8267

module ADD_8267 (
  input      [49:0]   io_A_0,
  input      [49:0]   io_A_1,
  input               io_CIN,
  output     [50:0]   io_S
);

  wire       [50:0]   _zz_io_S;
  wire       [50:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {50'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//KaratsubaCore_1427 replaced by KaratsubaCore_1435

module KaratsubaCore_1426 (
  input      [50:0]   io_a_0,
  input      [50:0]   io_b_0,
  output     [101:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [101:0]  basic_mul_io_p;

  BasicMUL48_958 basic_mul (
    .io_a   (io_a_0[50:0]         ), //i
    .io_b   (io_b_0[50:0]         ), //i
    .io_p   (basic_mul_io_p[101:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign io_p = basic_mul_io_p;

endmodule

//KaratsubaCore_1425 replaced by KaratsubaCore_1435

//BADD_2814 replaced by BADD_2818

//BADD_2813 replaced by BADD_2820

//BADD_2812 replaced by BADD_2819

//BADD_2811 replaced by BADD_2818

//ADD_8270 replaced by ADD_8288

//ADD_8269 replaced by ADD_8288

//KaratsubaCore_1430 replaced by KaratsubaCore_1438

//KaratsubaCore_1429 replaced by KaratsubaCore_1435

//KaratsubaCore_1428 replaced by KaratsubaCore_1438

//ADD_8276 replaced by ADD_11602

//ADD_8275 replaced by ADD_11602

//ADD_8274 replaced by ADD_11602

//ADD_8273 replaced by ADD_11602

//ADD_8272 replaced by ADD_11602

//ADD_8271 replaced by ADD_11602

//ADD_8281 replaced by ADD_11601

//ADD_8280 replaced by ADD_11602

//ADD_8279 replaced by ADD_11602

//ADD_8278 replaced by ADD_11602

//ADD_8277 replaced by ADD_11602

//ADD_8285 replaced by ADD_11602

//ADD_8284 replaced by ADD_11602

//ADD_8283 replaced by ADD_11602

//ADD_8282 replaced by ADD_11602

//BADD_2817 replaced by BADD_2824

//BADD_2816 replaced by BADD_2823

//BADD_2815 replaced by BADD_2822

//ADD_8287 replaced by ADD_11602

//ADD_8286 replaced by ADD_11602

//KaratsubaCore_1433 replaced by KaratsubaCore_1437

//KaratsubaCore_1432 replaced by KaratsubaCore_1438

//KaratsubaCore_1431 replaced by KaratsubaCore_1437

//BADD_2821 replaced by BADD_2818

module BADD_2820 (
  input      [98:0]   io_a,
  input      [98:0]   io_b,
  input               io_c,
  output     [99:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [2:0]    adder_adds_2_io_A_0;
  wire       [2:0]    adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [3:0]    adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [2:0]    _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11592 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[2:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[2:0]), //i
    .io_CIN (_zz_io_CIN_1            ), //i
    .io_S   (adder_adds_2_io_S[3:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[98 : 96];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[98 : 96];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_s <= adder_adds_2_io_S[3];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[2 : 0];
  end


endmodule

module BADD_2819 (
  input      [98:0]   io_a,
  input      [98:0]   io_b,
  input               io_c,
  output     [99:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [2:0]    adder_adds_2_io_A_0;
  wire       [2:0]    adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [3:0]    adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [2:0]    _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11592 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[2:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[2:0]), //i
    .io_CIN (_zz_io_CIN_1            ), //i
    .io_S   (adder_adds_2_io_S[3:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[98 : 96];
  assign adder_adds_0_io_A_1 = (~ io_b[47 : 0]);
  assign adder_adds_1_io_A_1 = (~ io_b[95 : 48]);
  assign adder_adds_2_io_A_1 = (~ io_b[98 : 96]);
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_s <= (! adder_adds_2_io_S[3]);
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[2 : 0];
  end


endmodule

module BADD_2818 (
  input      [97:0]   io_a,
  input      [97:0]   io_b,
  input               io_c,
  output     [98:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [1:0]    adder_adds_2_io_A_0;
  wire       [1:0]    adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [2:0]    adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [1:0]    _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11595 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[1:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[1:0]), //i
    .io_CIN (_zz_io_CIN_1            ), //i
    .io_S   (adder_adds_2_io_S[2:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[97 : 96];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[97 : 96];
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_s <= adder_adds_2_io_S[2];
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[1 : 0];
  end


endmodule

//ADD_8289 replaced by ADD_8288

module ADD_8288 (
  input      [48:0]   io_A_0,
  input      [48:0]   io_A_1,
  input               io_CIN,
  output     [49:0]   io_S
);

  wire       [49:0]   _zz_io_S;
  wire       [49:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {49'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//KaratsubaCore_1436 replaced by KaratsubaCore_1438

module KaratsubaCore_1435 (
  input      [49:0]   io_a_0,
  input      [49:0]   io_b_0,
  output     [99:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [99:0]   basic_mul_io_p;

  BasicMUL48_967 basic_mul (
    .io_a   (io_a_0[49:0]        ), //i
    .io_b   (io_b_0[49:0]        ), //i
    .io_p   (basic_mul_io_p[99:0]), //o
    .clk    (clk                 ), //i
    .resetn (resetn              )  //i
  );
  assign io_p = basic_mul_io_p;

endmodule

//KaratsubaCore_1434 replaced by KaratsubaCore_1438

module BADD_2824 (
  input      [143:0]  io_a,
  input      [143:0]  io_b,
  input               io_c,
  output     [144:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [47:0]   adder_adds_2_io_A_0;
  wire       [47:0]   adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [48:0]   adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg                 _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_2_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN_1             ), //i
    .io_S   (adder_adds_2_io_S[48:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[143 : 96];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign adder_adds_2_io_A_1 = io_b[143 : 96];
  assign io_s = {_zz_io_s_1,{_zz_io_s_4,{_zz_io_s_3,_zz_io_s_2}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_s <= adder_adds_2_io_S[48];
    _zz_io_s_1 <= _zz_io_s;
    _zz_io_s_2 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_4 <= adder_adds_2_io_S[47 : 0];
  end


endmodule

module BADD_2823 (
  input      [96:0]   io_a,
  input      [96:0]   io_b,
  input               io_c,
  output     [97:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [0:0]    adder_adds_2_io_A_0;
  wire       [0:0]    adder_adds_2_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  wire       [1:0]    adder_adds_2_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_CIN_1;
  reg                 _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [0:0]    _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  ADD_11601 adder_adds_2 (
    .io_A_0 (adder_adds_2_io_A_0   ), //i
    .io_A_1 (adder_adds_2_io_A_1   ), //i
    .io_CIN (_zz_io_CIN_1          ), //i
    .io_S   (adder_adds_2_io_S[1:0])  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_2_io_A_0 = io_a[96 : 96];
  assign adder_adds_0_io_A_1 = (~ io_b[47 : 0]);
  assign adder_adds_1_io_A_1 = (~ io_b[95 : 48]);
  assign adder_adds_2_io_A_1 = (~ io_b[96 : 96]);
  assign io_s = {_zz_io_s,{_zz_io_s_3,{_zz_io_s_2,_zz_io_s_1}}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_CIN_1 <= adder_adds_1_io_S[48];
    _zz_io_s <= (! adder_adds_2_io_S[1]);
    _zz_io_s_1 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_2 <= adder_adds_1_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_2_io_S[0 : 0];
  end


endmodule

module BADD_2822 (
  input      [95:0]   io_a,
  input      [95:0]   io_b,
  input               io_c,
  output     [96:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   adder_adds_0_io_A_0;
  wire       [47:0]   adder_adds_0_io_A_1;
  wire       [47:0]   adder_adds_1_io_A_0;
  wire       [47:0]   adder_adds_1_io_A_1;
  wire       [48:0]   adder_adds_0_io_S;
  wire       [48:0]   adder_adds_1_io_S;
  reg                 _zz_io_CIN;
  reg                 _zz_io_s;
  reg                 _zz_io_s_1;
  reg        [47:0]   _zz_io_s_2;
  reg        [47:0]   _zz_io_s_3;

  ADD_11602 adder_adds_0 (
    .io_A_0 (adder_adds_0_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_0_io_A_1[47:0]), //i
    .io_CIN (io_c                     ), //i
    .io_S   (adder_adds_0_io_S[48:0]  )  //o
  );
  ADD_11602 adder_adds_1 (
    .io_A_0 (adder_adds_1_io_A_0[47:0]), //i
    .io_A_1 (adder_adds_1_io_A_1[47:0]), //i
    .io_CIN (_zz_io_CIN               ), //i
    .io_S   (adder_adds_1_io_S[48:0]  )  //o
  );
  assign adder_adds_0_io_A_0 = io_a[47 : 0];
  assign adder_adds_1_io_A_0 = io_a[95 : 48];
  assign adder_adds_0_io_A_1 = io_b[47 : 0];
  assign adder_adds_1_io_A_1 = io_b[95 : 48];
  assign io_s = {_zz_io_s_1,{_zz_io_s_3,_zz_io_s_2}};
  always @(posedge clk) begin
    _zz_io_CIN <= adder_adds_0_io_S[48];
    _zz_io_s <= adder_adds_1_io_S[48];
    _zz_io_s_1 <= _zz_io_s;
    _zz_io_s_2 <= adder_adds_0_io_S[47 : 0];
    _zz_io_s_3 <= adder_adds_1_io_S[47 : 0];
  end


endmodule

//ADD_8291 replaced by ADD_11602

//ADD_8290 replaced by ADD_11602

//KaratsubaCore_1439 replaced by KaratsubaCore_1437

module KaratsubaCore_1438 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_b_0,
  output     [97:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [97:0]   basic_mul_io_p;

  BasicMUL48_970 basic_mul (
    .io_a   (io_a_0[48:0]        ), //i
    .io_b   (io_b_0[48:0]        ), //i
    .io_p   (basic_mul_io_p[97:0]), //o
    .clk    (clk                 ), //i
    .resetn (resetn              )  //i
  );
  assign io_p = basic_mul_io_p;

endmodule

module KaratsubaCore_1437 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_b_0,
  output     [95:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [95:0]   basic_mul_io_p;

  BasicMUL48_971 basic_mul (
    .io_a   (io_a_0[47:0]        ), //i
    .io_b   (io_b_0[47:0]        ), //i
    .io_p   (basic_mul_io_p[95:0]), //o
    .clk    (clk                 ), //i
    .resetn (resetn              )  //i
  );
  assign io_p = basic_mul_io_p;

endmodule

//ADD_8294 replaced by ADD_11602

//ADD_8293 replaced by ADD_11602

//ADD_8292 replaced by ADD_11602

//ADD_8297 replaced by ADD_11601

//ADD_8296 replaced by ADD_11602

//ADD_8295 replaced by ADD_11602

//ADD_8299 replaced by ADD_11602

//ADD_8298 replaced by ADD_11602

//BasicMUL48 replaced by BasicMUL48_971

//BasicMUL48_1 replaced by BasicMUL48_970

//BasicMUL48_2 replaced by BasicMUL48_971

//ADD_8302 replaced by ADD_11595

//ADD_8301 replaced by ADD_11602

//ADD_8300 replaced by ADD_11602

//ADD_8305 replaced by ADD_11592

//ADD_8304 replaced by ADD_11602

//ADD_8303 replaced by ADD_11602

//ADD_8308 replaced by ADD_11592

//ADD_8307 replaced by ADD_11602

//ADD_8306 replaced by ADD_11602

//ADD_8311 replaced by ADD_11595

//ADD_8310 replaced by ADD_11602

//ADD_8309 replaced by ADD_11602

//BasicMUL48_3 replaced by BasicMUL48_970

//BasicMUL48_4 replaced by BasicMUL48_967

//BasicMUL48_5 replaced by BasicMUL48_970

//ADD_8314 replaced by ADD_11602

//ADD_8313 replaced by ADD_11602

//ADD_8312 replaced by ADD_11602

//ADD_8317 replaced by ADD_11601

//ADD_8316 replaced by ADD_11602

//ADD_8315 replaced by ADD_11602

//ADD_8319 replaced by ADD_11602

//ADD_8318 replaced by ADD_11602

//BasicMUL48_6 replaced by BasicMUL48_971

//BasicMUL48_7 replaced by BasicMUL48_970

//BasicMUL48_8 replaced by BasicMUL48_971

//ADD_8322 replaced by ADD_11595

//ADD_8321 replaced by ADD_11602

//ADD_8320 replaced by ADD_11602

//ADD_8325 replaced by ADD_11592

//ADD_8324 replaced by ADD_11602

//ADD_8323 replaced by ADD_11602

//ADD_8328 replaced by ADD_11592

//ADD_8327 replaced by ADD_11602

//ADD_8326 replaced by ADD_11602

//ADD_8331 replaced by ADD_11595

//ADD_8330 replaced by ADD_11602

//ADD_8329 replaced by ADD_11602

//BasicMUL48_9 replaced by BasicMUL48_970

//BasicMUL48_10 replaced by BasicMUL48_967

//BasicMUL48_11 replaced by BasicMUL48_970

//ADD_8334 replaced by ADD_11563

//ADD_8333 replaced by ADD_11602

//ADD_8332 replaced by ADD_11602

//ADD_8337 replaced by ADD_11560

//ADD_8336 replaced by ADD_11602

//ADD_8335 replaced by ADD_11602

//ADD_8340 replaced by ADD_11560

//ADD_8339 replaced by ADD_11602

//ADD_8338 replaced by ADD_11602

//ADD_8343 replaced by ADD_11563

//ADD_8342 replaced by ADD_11602

//ADD_8341 replaced by ADD_11602

//BasicMUL48_12 replaced by BasicMUL48_967

//BasicMUL48_13 replaced by BasicMUL48_958

//BasicMUL48_14 replaced by BasicMUL48_967

//ADD_8346 replaced by ADD_11595

//ADD_8345 replaced by ADD_11602

//ADD_8344 replaced by ADD_11602

//ADD_8349 replaced by ADD_11592

//ADD_8348 replaced by ADD_11602

//ADD_8347 replaced by ADD_11602

//ADD_8352 replaced by ADD_11592

//ADD_8351 replaced by ADD_11602

//ADD_8350 replaced by ADD_11602

//ADD_8355 replaced by ADD_11595

//ADD_8354 replaced by ADD_11602

//ADD_8353 replaced by ADD_11602

//BasicMUL48_15 replaced by BasicMUL48_970

//BasicMUL48_16 replaced by BasicMUL48_967

//BasicMUL48_17 replaced by BasicMUL48_970

//ADD_8358 replaced by ADD_11602

//ADD_8357 replaced by ADD_11602

//ADD_8356 replaced by ADD_11602

//ADD_8361 replaced by ADD_11601

//ADD_8360 replaced by ADD_11602

//ADD_8359 replaced by ADD_11602

//ADD_8363 replaced by ADD_11602

//ADD_8362 replaced by ADD_11602

//BasicMUL48_18 replaced by BasicMUL48_971

//BasicMUL48_19 replaced by BasicMUL48_970

//BasicMUL48_20 replaced by BasicMUL48_971

//ADD_8366 replaced by ADD_11595

//ADD_8365 replaced by ADD_11602

//ADD_8364 replaced by ADD_11602

//ADD_8369 replaced by ADD_11592

//ADD_8368 replaced by ADD_11602

//ADD_8367 replaced by ADD_11602

//ADD_8372 replaced by ADD_11592

//ADD_8371 replaced by ADD_11602

//ADD_8370 replaced by ADD_11602

//ADD_8375 replaced by ADD_11595

//ADD_8374 replaced by ADD_11602

//ADD_8373 replaced by ADD_11602

//BasicMUL48_21 replaced by BasicMUL48_970

//BasicMUL48_22 replaced by BasicMUL48_967

//BasicMUL48_23 replaced by BasicMUL48_970

//ADD_8378 replaced by ADD_11602

//ADD_8377 replaced by ADD_11602

//ADD_8376 replaced by ADD_11602

//ADD_8381 replaced by ADD_11601

//ADD_8380 replaced by ADD_11602

//ADD_8379 replaced by ADD_11602

//ADD_8383 replaced by ADD_11602

//ADD_8382 replaced by ADD_11602

//BasicMUL48_24 replaced by BasicMUL48_971

//BasicMUL48_25 replaced by BasicMUL48_970

//BasicMUL48_26 replaced by BasicMUL48_971

//ADD_8386 replaced by ADD_11602

//ADD_8385 replaced by ADD_11602

//ADD_8384 replaced by ADD_11602

//ADD_8389 replaced by ADD_11601

//ADD_8388 replaced by ADD_11602

//ADD_8387 replaced by ADD_11602

//ADD_8391 replaced by ADD_11602

//ADD_8390 replaced by ADD_11602

//BasicMUL48_27 replaced by BasicMUL48_971

//BasicMUL48_28 replaced by BasicMUL48_970

//BasicMUL48_29 replaced by BasicMUL48_971

//ADD_8394 replaced by ADD_11595

//ADD_8393 replaced by ADD_11602

//ADD_8392 replaced by ADD_11602

//ADD_8397 replaced by ADD_11592

//ADD_8396 replaced by ADD_11602

//ADD_8395 replaced by ADD_11602

//ADD_8400 replaced by ADD_11592

//ADD_8399 replaced by ADD_11602

//ADD_8398 replaced by ADD_11602

//ADD_8403 replaced by ADD_11595

//ADD_8402 replaced by ADD_11602

//ADD_8401 replaced by ADD_11602

//BasicMUL48_30 replaced by BasicMUL48_970

//BasicMUL48_31 replaced by BasicMUL48_967

//BasicMUL48_32 replaced by BasicMUL48_970

//ADD_8406 replaced by ADD_11602

//ADD_8405 replaced by ADD_11602

//ADD_8404 replaced by ADD_11602

//ADD_8409 replaced by ADD_11601

//ADD_8408 replaced by ADD_11602

//ADD_8407 replaced by ADD_11602

//ADD_8411 replaced by ADD_11602

//ADD_8410 replaced by ADD_11602

//BasicMUL48_33 replaced by BasicMUL48_971

//BasicMUL48_34 replaced by BasicMUL48_970

//BasicMUL48_35 replaced by BasicMUL48_971

//ADD_8414 replaced by ADD_11595

//ADD_8413 replaced by ADD_11602

//ADD_8412 replaced by ADD_11602

//ADD_8417 replaced by ADD_11592

//ADD_8416 replaced by ADD_11602

//ADD_8415 replaced by ADD_11602

//ADD_8420 replaced by ADD_11592

//ADD_8419 replaced by ADD_11602

//ADD_8418 replaced by ADD_11602

//ADD_8423 replaced by ADD_11595

//ADD_8422 replaced by ADD_11602

//ADD_8421 replaced by ADD_11602

//BasicMUL48_36 replaced by BasicMUL48_970

//BasicMUL48_37 replaced by BasicMUL48_967

//BasicMUL48_38 replaced by BasicMUL48_970

//ADD_8426 replaced by ADD_11563

//ADD_8425 replaced by ADD_11602

//ADD_8424 replaced by ADD_11602

//ADD_8429 replaced by ADD_11560

//ADD_8428 replaced by ADD_11602

//ADD_8427 replaced by ADD_11602

//ADD_8432 replaced by ADD_11560

//ADD_8431 replaced by ADD_11602

//ADD_8430 replaced by ADD_11602

//ADD_8435 replaced by ADD_11563

//ADD_8434 replaced by ADD_11602

//ADD_8433 replaced by ADD_11602

//BasicMUL48_39 replaced by BasicMUL48_967

//BasicMUL48_40 replaced by BasicMUL48_958

//BasicMUL48_41 replaced by BasicMUL48_967

//ADD_8438 replaced by ADD_11595

//ADD_8437 replaced by ADD_11602

//ADD_8436 replaced by ADD_11602

//ADD_8441 replaced by ADD_11592

//ADD_8440 replaced by ADD_11602

//ADD_8439 replaced by ADD_11602

//ADD_8444 replaced by ADD_11592

//ADD_8443 replaced by ADD_11602

//ADD_8442 replaced by ADD_11602

//ADD_8447 replaced by ADD_11595

//ADD_8446 replaced by ADD_11602

//ADD_8445 replaced by ADD_11602

//BasicMUL48_42 replaced by BasicMUL48_970

//BasicMUL48_43 replaced by BasicMUL48_967

//BasicMUL48_44 replaced by BasicMUL48_970

//ADD_8450 replaced by ADD_11602

//ADD_8449 replaced by ADD_11602

//ADD_8448 replaced by ADD_11602

//ADD_8453 replaced by ADD_11601

//ADD_8452 replaced by ADD_11602

//ADD_8451 replaced by ADD_11602

//ADD_8455 replaced by ADD_11602

//ADD_8454 replaced by ADD_11602

//BasicMUL48_45 replaced by BasicMUL48_971

//BasicMUL48_46 replaced by BasicMUL48_970

//BasicMUL48_47 replaced by BasicMUL48_971

//ADD_8458 replaced by ADD_11595

//ADD_8457 replaced by ADD_11602

//ADD_8456 replaced by ADD_11602

//ADD_8461 replaced by ADD_11592

//ADD_8460 replaced by ADD_11602

//ADD_8459 replaced by ADD_11602

//ADD_8464 replaced by ADD_11592

//ADD_8463 replaced by ADD_11602

//ADD_8462 replaced by ADD_11602

//ADD_8467 replaced by ADD_11595

//ADD_8466 replaced by ADD_11602

//ADD_8465 replaced by ADD_11602

//BasicMUL48_48 replaced by BasicMUL48_970

//BasicMUL48_49 replaced by BasicMUL48_967

//BasicMUL48_50 replaced by BasicMUL48_970

//ADD_8470 replaced by ADD_11602

//ADD_8469 replaced by ADD_11602

//ADD_8468 replaced by ADD_11602

//ADD_8473 replaced by ADD_11601

//ADD_8472 replaced by ADD_11602

//ADD_8471 replaced by ADD_11602

//ADD_8475 replaced by ADD_11602

//ADD_8474 replaced by ADD_11602

//BasicMUL48_51 replaced by BasicMUL48_971

//BasicMUL48_52 replaced by BasicMUL48_970

//BasicMUL48_53 replaced by BasicMUL48_971

//ADD_8478 replaced by ADD_11602

//ADD_8477 replaced by ADD_11602

//ADD_8476 replaced by ADD_11602

//ADD_8481 replaced by ADD_11601

//ADD_8480 replaced by ADD_11602

//ADD_8479 replaced by ADD_11602

//ADD_8483 replaced by ADD_11602

//ADD_8482 replaced by ADD_11602

//BasicMUL48_54 replaced by BasicMUL48_971

//BasicMUL48_55 replaced by BasicMUL48_970

//BasicMUL48_56 replaced by BasicMUL48_971

//ADD_8486 replaced by ADD_11595

//ADD_8485 replaced by ADD_11602

//ADD_8484 replaced by ADD_11602

//ADD_8489 replaced by ADD_11592

//ADD_8488 replaced by ADD_11602

//ADD_8487 replaced by ADD_11602

//ADD_8492 replaced by ADD_11592

//ADD_8491 replaced by ADD_11602

//ADD_8490 replaced by ADD_11602

//ADD_8495 replaced by ADD_11595

//ADD_8494 replaced by ADD_11602

//ADD_8493 replaced by ADD_11602

//BasicMUL48_57 replaced by BasicMUL48_970

//BasicMUL48_58 replaced by BasicMUL48_967

//BasicMUL48_59 replaced by BasicMUL48_970

//ADD_8498 replaced by ADD_11602

//ADD_8497 replaced by ADD_11602

//ADD_8496 replaced by ADD_11602

//ADD_8501 replaced by ADD_11601

//ADD_8500 replaced by ADD_11602

//ADD_8499 replaced by ADD_11602

//ADD_8503 replaced by ADD_11602

//ADD_8502 replaced by ADD_11602

//BasicMUL48_60 replaced by BasicMUL48_971

//BasicMUL48_61 replaced by BasicMUL48_970

//BasicMUL48_62 replaced by BasicMUL48_971

//ADD_8506 replaced by ADD_11595

//ADD_8505 replaced by ADD_11602

//ADD_8504 replaced by ADD_11602

//ADD_8509 replaced by ADD_11592

//ADD_8508 replaced by ADD_11602

//ADD_8507 replaced by ADD_11602

//ADD_8512 replaced by ADD_11592

//ADD_8511 replaced by ADD_11602

//ADD_8510 replaced by ADD_11602

//ADD_8515 replaced by ADD_11595

//ADD_8514 replaced by ADD_11602

//ADD_8513 replaced by ADD_11602

//BasicMUL48_63 replaced by BasicMUL48_970

//BasicMUL48_64 replaced by BasicMUL48_967

//BasicMUL48_65 replaced by BasicMUL48_970

//ADD_8518 replaced by ADD_11563

//ADD_8517 replaced by ADD_11602

//ADD_8516 replaced by ADD_11602

//ADD_8521 replaced by ADD_11560

//ADD_8520 replaced by ADD_11602

//ADD_8519 replaced by ADD_11602

//ADD_8524 replaced by ADD_11560

//ADD_8523 replaced by ADD_11602

//ADD_8522 replaced by ADD_11602

//ADD_8527 replaced by ADD_11563

//ADD_8526 replaced by ADD_11602

//ADD_8525 replaced by ADD_11602

//BasicMUL48_66 replaced by BasicMUL48_967

//BasicMUL48_67 replaced by BasicMUL48_958

//BasicMUL48_68 replaced by BasicMUL48_967

//ADD_8530 replaced by ADD_11595

//ADD_8529 replaced by ADD_11602

//ADD_8528 replaced by ADD_11602

//ADD_8533 replaced by ADD_11592

//ADD_8532 replaced by ADD_11602

//ADD_8531 replaced by ADD_11602

//ADD_8536 replaced by ADD_11592

//ADD_8535 replaced by ADD_11602

//ADD_8534 replaced by ADD_11602

//ADD_8539 replaced by ADD_11595

//ADD_8538 replaced by ADD_11602

//ADD_8537 replaced by ADD_11602

//BasicMUL48_69 replaced by BasicMUL48_970

//BasicMUL48_70 replaced by BasicMUL48_967

//BasicMUL48_71 replaced by BasicMUL48_970

//ADD_8542 replaced by ADD_11602

//ADD_8541 replaced by ADD_11602

//ADD_8540 replaced by ADD_11602

//ADD_8545 replaced by ADD_11601

//ADD_8544 replaced by ADD_11602

//ADD_8543 replaced by ADD_11602

//ADD_8547 replaced by ADD_11602

//ADD_8546 replaced by ADD_11602

//BasicMUL48_72 replaced by BasicMUL48_971

//BasicMUL48_73 replaced by BasicMUL48_970

//BasicMUL48_74 replaced by BasicMUL48_971

//ADD_8550 replaced by ADD_11595

//ADD_8549 replaced by ADD_11602

//ADD_8548 replaced by ADD_11602

//ADD_8553 replaced by ADD_11592

//ADD_8552 replaced by ADD_11602

//ADD_8551 replaced by ADD_11602

//ADD_8556 replaced by ADD_11592

//ADD_8555 replaced by ADD_11602

//ADD_8554 replaced by ADD_11602

//ADD_8559 replaced by ADD_11595

//ADD_8558 replaced by ADD_11602

//ADD_8557 replaced by ADD_11602

//BasicMUL48_75 replaced by BasicMUL48_970

//BasicMUL48_76 replaced by BasicMUL48_967

//BasicMUL48_77 replaced by BasicMUL48_970

//ADD_8562 replaced by ADD_11602

//ADD_8561 replaced by ADD_11602

//ADD_8560 replaced by ADD_11602

//ADD_8565 replaced by ADD_11601

//ADD_8564 replaced by ADD_11602

//ADD_8563 replaced by ADD_11602

//ADD_8567 replaced by ADD_11602

//ADD_8566 replaced by ADD_11602

//BasicMUL48_78 replaced by BasicMUL48_971

//BasicMUL48_79 replaced by BasicMUL48_970

//BasicMUL48_80 replaced by BasicMUL48_971

//ADD_8570 replaced by ADD_11602

//ADD_8569 replaced by ADD_11602

//ADD_8568 replaced by ADD_11602

//ADD_8573 replaced by ADD_11601

//ADD_8572 replaced by ADD_11602

//ADD_8571 replaced by ADD_11602

//ADD_8575 replaced by ADD_11602

//ADD_8574 replaced by ADD_11602

//BasicMUL48_81 replaced by BasicMUL48_971

//BasicMUL48_82 replaced by BasicMUL48_970

//BasicMUL48_83 replaced by BasicMUL48_971

//ADD_8578 replaced by ADD_11595

//ADD_8577 replaced by ADD_11602

//ADD_8576 replaced by ADD_11602

//ADD_8581 replaced by ADD_11592

//ADD_8580 replaced by ADD_11602

//ADD_8579 replaced by ADD_11602

//ADD_8584 replaced by ADD_11592

//ADD_8583 replaced by ADD_11602

//ADD_8582 replaced by ADD_11602

//ADD_8587 replaced by ADD_11595

//ADD_8586 replaced by ADD_11602

//ADD_8585 replaced by ADD_11602

//BasicMUL48_84 replaced by BasicMUL48_970

//BasicMUL48_85 replaced by BasicMUL48_967

//BasicMUL48_86 replaced by BasicMUL48_970

//ADD_8590 replaced by ADD_11602

//ADD_8589 replaced by ADD_11602

//ADD_8588 replaced by ADD_11602

//ADD_8593 replaced by ADD_11601

//ADD_8592 replaced by ADD_11602

//ADD_8591 replaced by ADD_11602

//ADD_8595 replaced by ADD_11602

//ADD_8594 replaced by ADD_11602

//BasicMUL48_87 replaced by BasicMUL48_971

//BasicMUL48_88 replaced by BasicMUL48_970

//BasicMUL48_89 replaced by BasicMUL48_971

//ADD_8598 replaced by ADD_11595

//ADD_8597 replaced by ADD_11602

//ADD_8596 replaced by ADD_11602

//ADD_8601 replaced by ADD_11592

//ADD_8600 replaced by ADD_11602

//ADD_8599 replaced by ADD_11602

//ADD_8604 replaced by ADD_11592

//ADD_8603 replaced by ADD_11602

//ADD_8602 replaced by ADD_11602

//ADD_8607 replaced by ADD_11595

//ADD_8606 replaced by ADD_11602

//ADD_8605 replaced by ADD_11602

//BasicMUL48_90 replaced by BasicMUL48_970

//BasicMUL48_91 replaced by BasicMUL48_967

//BasicMUL48_92 replaced by BasicMUL48_970

//ADD_8610 replaced by ADD_11563

//ADD_8609 replaced by ADD_11602

//ADD_8608 replaced by ADD_11602

//ADD_8613 replaced by ADD_11560

//ADD_8612 replaced by ADD_11602

//ADD_8611 replaced by ADD_11602

//ADD_8616 replaced by ADD_11560

//ADD_8615 replaced by ADD_11602

//ADD_8614 replaced by ADD_11602

//ADD_8619 replaced by ADD_11563

//ADD_8618 replaced by ADD_11602

//ADD_8617 replaced by ADD_11602

//BasicMUL48_93 replaced by BasicMUL48_967

//BasicMUL48_94 replaced by BasicMUL48_958

//BasicMUL48_95 replaced by BasicMUL48_967

//ADD_8622 replaced by ADD_11595

//ADD_8621 replaced by ADD_11602

//ADD_8620 replaced by ADD_11602

//ADD_8625 replaced by ADD_11592

//ADD_8624 replaced by ADD_11602

//ADD_8623 replaced by ADD_11602

//ADD_8628 replaced by ADD_11592

//ADD_8627 replaced by ADD_11602

//ADD_8626 replaced by ADD_11602

//ADD_8631 replaced by ADD_11595

//ADD_8630 replaced by ADD_11602

//ADD_8629 replaced by ADD_11602

//BasicMUL48_96 replaced by BasicMUL48_970

//BasicMUL48_97 replaced by BasicMUL48_967

//BasicMUL48_98 replaced by BasicMUL48_970

//ADD_8634 replaced by ADD_11602

//ADD_8633 replaced by ADD_11602

//ADD_8632 replaced by ADD_11602

//ADD_8637 replaced by ADD_11601

//ADD_8636 replaced by ADD_11602

//ADD_8635 replaced by ADD_11602

//ADD_8639 replaced by ADD_11602

//ADD_8638 replaced by ADD_11602

//BasicMUL48_99 replaced by BasicMUL48_971

//BasicMUL48_100 replaced by BasicMUL48_970

//BasicMUL48_101 replaced by BasicMUL48_971

//ADD_8642 replaced by ADD_11595

//ADD_8641 replaced by ADD_11602

//ADD_8640 replaced by ADD_11602

//ADD_8645 replaced by ADD_11592

//ADD_8644 replaced by ADD_11602

//ADD_8643 replaced by ADD_11602

//ADD_8648 replaced by ADD_11592

//ADD_8647 replaced by ADD_11602

//ADD_8646 replaced by ADD_11602

//ADD_8651 replaced by ADD_11595

//ADD_8650 replaced by ADD_11602

//ADD_8649 replaced by ADD_11602

//BasicMUL48_102 replaced by BasicMUL48_970

//BasicMUL48_103 replaced by BasicMUL48_967

//BasicMUL48_104 replaced by BasicMUL48_970

//ADD_8654 replaced by ADD_11602

//ADD_8653 replaced by ADD_11602

//ADD_8652 replaced by ADD_11602

//ADD_8657 replaced by ADD_11601

//ADD_8656 replaced by ADD_11602

//ADD_8655 replaced by ADD_11602

//ADD_8659 replaced by ADD_11602

//ADD_8658 replaced by ADD_11602

//BasicMUL48_105 replaced by BasicMUL48_971

//BasicMUL48_106 replaced by BasicMUL48_970

//BasicMUL48_107 replaced by BasicMUL48_971

//ADD_8662 replaced by ADD_11602

//ADD_8661 replaced by ADD_11602

//ADD_8660 replaced by ADD_11602

//ADD_8665 replaced by ADD_11601

//ADD_8664 replaced by ADD_11602

//ADD_8663 replaced by ADD_11602

//ADD_8667 replaced by ADD_11602

//ADD_8666 replaced by ADD_11602

//BasicMUL48_108 replaced by BasicMUL48_971

//BasicMUL48_109 replaced by BasicMUL48_970

//BasicMUL48_110 replaced by BasicMUL48_971

//ADD_8670 replaced by ADD_11595

//ADD_8669 replaced by ADD_11602

//ADD_8668 replaced by ADD_11602

//ADD_8673 replaced by ADD_11592

//ADD_8672 replaced by ADD_11602

//ADD_8671 replaced by ADD_11602

//ADD_8676 replaced by ADD_11592

//ADD_8675 replaced by ADD_11602

//ADD_8674 replaced by ADD_11602

//ADD_8679 replaced by ADD_11595

//ADD_8678 replaced by ADD_11602

//ADD_8677 replaced by ADD_11602

//BasicMUL48_111 replaced by BasicMUL48_970

//BasicMUL48_112 replaced by BasicMUL48_967

//BasicMUL48_113 replaced by BasicMUL48_970

//ADD_8682 replaced by ADD_11602

//ADD_8681 replaced by ADD_11602

//ADD_8680 replaced by ADD_11602

//ADD_8685 replaced by ADD_11601

//ADD_8684 replaced by ADD_11602

//ADD_8683 replaced by ADD_11602

//ADD_8687 replaced by ADD_11602

//ADD_8686 replaced by ADD_11602

//BasicMUL48_114 replaced by BasicMUL48_971

//BasicMUL48_115 replaced by BasicMUL48_970

//BasicMUL48_116 replaced by BasicMUL48_971

//ADD_8690 replaced by ADD_11595

//ADD_8689 replaced by ADD_11602

//ADD_8688 replaced by ADD_11602

//ADD_8693 replaced by ADD_11592

//ADD_8692 replaced by ADD_11602

//ADD_8691 replaced by ADD_11602

//ADD_8696 replaced by ADD_11592

//ADD_8695 replaced by ADD_11602

//ADD_8694 replaced by ADD_11602

//ADD_8699 replaced by ADD_11595

//ADD_8698 replaced by ADD_11602

//ADD_8697 replaced by ADD_11602

//BasicMUL48_117 replaced by BasicMUL48_970

//BasicMUL48_118 replaced by BasicMUL48_967

//BasicMUL48_119 replaced by BasicMUL48_970

//ADD_8702 replaced by ADD_11563

//ADD_8701 replaced by ADD_11602

//ADD_8700 replaced by ADD_11602

//ADD_8705 replaced by ADD_11560

//ADD_8704 replaced by ADD_11602

//ADD_8703 replaced by ADD_11602

//ADD_8708 replaced by ADD_11560

//ADD_8707 replaced by ADD_11602

//ADD_8706 replaced by ADD_11602

//ADD_8711 replaced by ADD_11563

//ADD_8710 replaced by ADD_11602

//ADD_8709 replaced by ADD_11602

//BasicMUL48_120 replaced by BasicMUL48_967

//BasicMUL48_121 replaced by BasicMUL48_958

//BasicMUL48_122 replaced by BasicMUL48_967

//ADD_8714 replaced by ADD_11595

//ADD_8713 replaced by ADD_11602

//ADD_8712 replaced by ADD_11602

//ADD_8717 replaced by ADD_11592

//ADD_8716 replaced by ADD_11602

//ADD_8715 replaced by ADD_11602

//ADD_8720 replaced by ADD_11592

//ADD_8719 replaced by ADD_11602

//ADD_8718 replaced by ADD_11602

//ADD_8723 replaced by ADD_11595

//ADD_8722 replaced by ADD_11602

//ADD_8721 replaced by ADD_11602

//BasicMUL48_123 replaced by BasicMUL48_970

//BasicMUL48_124 replaced by BasicMUL48_967

//BasicMUL48_125 replaced by BasicMUL48_970

//ADD_8726 replaced by ADD_11602

//ADD_8725 replaced by ADD_11602

//ADD_8724 replaced by ADD_11602

//ADD_8729 replaced by ADD_11601

//ADD_8728 replaced by ADD_11602

//ADD_8727 replaced by ADD_11602

//ADD_8731 replaced by ADD_11602

//ADD_8730 replaced by ADD_11602

//BasicMUL48_126 replaced by BasicMUL48_971

//BasicMUL48_127 replaced by BasicMUL48_970

//BasicMUL48_128 replaced by BasicMUL48_971

//ADD_8734 replaced by ADD_11595

//ADD_8733 replaced by ADD_11602

//ADD_8732 replaced by ADD_11602

//ADD_8737 replaced by ADD_11592

//ADD_8736 replaced by ADD_11602

//ADD_8735 replaced by ADD_11602

//ADD_8740 replaced by ADD_11592

//ADD_8739 replaced by ADD_11602

//ADD_8738 replaced by ADD_11602

//ADD_8743 replaced by ADD_11595

//ADD_8742 replaced by ADD_11602

//ADD_8741 replaced by ADD_11602

//BasicMUL48_129 replaced by BasicMUL48_970

//BasicMUL48_130 replaced by BasicMUL48_967

//BasicMUL48_131 replaced by BasicMUL48_970

//ADD_8746 replaced by ADD_11602

//ADD_8745 replaced by ADD_11602

//ADD_8744 replaced by ADD_11602

//ADD_8749 replaced by ADD_11601

//ADD_8748 replaced by ADD_11602

//ADD_8747 replaced by ADD_11602

//ADD_8751 replaced by ADD_11602

//ADD_8750 replaced by ADD_11602

//BasicMUL48_132 replaced by BasicMUL48_971

//BasicMUL48_133 replaced by BasicMUL48_970

//BasicMUL48_134 replaced by BasicMUL48_971

//ADD_8754 replaced by ADD_11602

//ADD_8753 replaced by ADD_11602

//ADD_8752 replaced by ADD_11602

//ADD_8757 replaced by ADD_11601

//ADD_8756 replaced by ADD_11602

//ADD_8755 replaced by ADD_11602

//ADD_8759 replaced by ADD_11602

//ADD_8758 replaced by ADD_11602

//BasicMUL48_135 replaced by BasicMUL48_971

//BasicMUL48_136 replaced by BasicMUL48_970

//BasicMUL48_137 replaced by BasicMUL48_971

//ADD_8762 replaced by ADD_11595

//ADD_8761 replaced by ADD_11602

//ADD_8760 replaced by ADD_11602

//ADD_8765 replaced by ADD_11592

//ADD_8764 replaced by ADD_11602

//ADD_8763 replaced by ADD_11602

//ADD_8768 replaced by ADD_11592

//ADD_8767 replaced by ADD_11602

//ADD_8766 replaced by ADD_11602

//ADD_8771 replaced by ADD_11595

//ADD_8770 replaced by ADD_11602

//ADD_8769 replaced by ADD_11602

//BasicMUL48_138 replaced by BasicMUL48_970

//BasicMUL48_139 replaced by BasicMUL48_967

//BasicMUL48_140 replaced by BasicMUL48_970

//ADD_8774 replaced by ADD_11602

//ADD_8773 replaced by ADD_11602

//ADD_8772 replaced by ADD_11602

//ADD_8777 replaced by ADD_11601

//ADD_8776 replaced by ADD_11602

//ADD_8775 replaced by ADD_11602

//ADD_8779 replaced by ADD_11602

//ADD_8778 replaced by ADD_11602

//BasicMUL48_141 replaced by BasicMUL48_971

//BasicMUL48_142 replaced by BasicMUL48_970

//BasicMUL48_143 replaced by BasicMUL48_971

//ADD_8782 replaced by ADD_11595

//ADD_8781 replaced by ADD_11602

//ADD_8780 replaced by ADD_11602

//ADD_8785 replaced by ADD_11592

//ADD_8784 replaced by ADD_11602

//ADD_8783 replaced by ADD_11602

//ADD_8788 replaced by ADD_11592

//ADD_8787 replaced by ADD_11602

//ADD_8786 replaced by ADD_11602

//ADD_8791 replaced by ADD_11595

//ADD_8790 replaced by ADD_11602

//ADD_8789 replaced by ADD_11602

//BasicMUL48_144 replaced by BasicMUL48_970

//BasicMUL48_145 replaced by BasicMUL48_967

//BasicMUL48_146 replaced by BasicMUL48_970

//ADD_8794 replaced by ADD_11563

//ADD_8793 replaced by ADD_11602

//ADD_8792 replaced by ADD_11602

//ADD_8797 replaced by ADD_11560

//ADD_8796 replaced by ADD_11602

//ADD_8795 replaced by ADD_11602

//ADD_8800 replaced by ADD_11560

//ADD_8799 replaced by ADD_11602

//ADD_8798 replaced by ADD_11602

//ADD_8803 replaced by ADD_11563

//ADD_8802 replaced by ADD_11602

//ADD_8801 replaced by ADD_11602

//BasicMUL48_147 replaced by BasicMUL48_967

//BasicMUL48_148 replaced by BasicMUL48_958

//BasicMUL48_149 replaced by BasicMUL48_967

//ADD_8806 replaced by ADD_11595

//ADD_8805 replaced by ADD_11602

//ADD_8804 replaced by ADD_11602

//ADD_8809 replaced by ADD_11592

//ADD_8808 replaced by ADD_11602

//ADD_8807 replaced by ADD_11602

//ADD_8812 replaced by ADD_11592

//ADD_8811 replaced by ADD_11602

//ADD_8810 replaced by ADD_11602

//ADD_8815 replaced by ADD_11595

//ADD_8814 replaced by ADD_11602

//ADD_8813 replaced by ADD_11602

//BasicMUL48_150 replaced by BasicMUL48_970

//BasicMUL48_151 replaced by BasicMUL48_967

//BasicMUL48_152 replaced by BasicMUL48_970

//ADD_8818 replaced by ADD_11602

//ADD_8817 replaced by ADD_11602

//ADD_8816 replaced by ADD_11602

//ADD_8821 replaced by ADD_11601

//ADD_8820 replaced by ADD_11602

//ADD_8819 replaced by ADD_11602

//ADD_8823 replaced by ADD_11602

//ADD_8822 replaced by ADD_11602

//BasicMUL48_153 replaced by BasicMUL48_971

//BasicMUL48_154 replaced by BasicMUL48_970

//BasicMUL48_155 replaced by BasicMUL48_971

//ADD_8826 replaced by ADD_11595

//ADD_8825 replaced by ADD_11602

//ADD_8824 replaced by ADD_11602

//ADD_8829 replaced by ADD_11592

//ADD_8828 replaced by ADD_11602

//ADD_8827 replaced by ADD_11602

//ADD_8832 replaced by ADD_11592

//ADD_8831 replaced by ADD_11602

//ADD_8830 replaced by ADD_11602

//ADD_8835 replaced by ADD_11595

//ADD_8834 replaced by ADD_11602

//ADD_8833 replaced by ADD_11602

//BasicMUL48_156 replaced by BasicMUL48_970

//BasicMUL48_157 replaced by BasicMUL48_967

//BasicMUL48_158 replaced by BasicMUL48_970

//ADD_8838 replaced by ADD_11602

//ADD_8837 replaced by ADD_11602

//ADD_8836 replaced by ADD_11602

//ADD_8841 replaced by ADD_11601

//ADD_8840 replaced by ADD_11602

//ADD_8839 replaced by ADD_11602

//ADD_8843 replaced by ADD_11602

//ADD_8842 replaced by ADD_11602

//BasicMUL48_159 replaced by BasicMUL48_971

//BasicMUL48_160 replaced by BasicMUL48_970

//BasicMUL48_161 replaced by BasicMUL48_971

//ADD_8846 replaced by ADD_11602

//ADD_8845 replaced by ADD_11602

//ADD_8844 replaced by ADD_11602

//ADD_8849 replaced by ADD_11601

//ADD_8848 replaced by ADD_11602

//ADD_8847 replaced by ADD_11602

//ADD_8851 replaced by ADD_11602

//ADD_8850 replaced by ADD_11602

//BasicMUL48_162 replaced by BasicMUL48_971

//BasicMUL48_163 replaced by BasicMUL48_970

//BasicMUL48_164 replaced by BasicMUL48_971

//ADD_8854 replaced by ADD_11595

//ADD_8853 replaced by ADD_11602

//ADD_8852 replaced by ADD_11602

//ADD_8857 replaced by ADD_11592

//ADD_8856 replaced by ADD_11602

//ADD_8855 replaced by ADD_11602

//ADD_8860 replaced by ADD_11592

//ADD_8859 replaced by ADD_11602

//ADD_8858 replaced by ADD_11602

//ADD_8863 replaced by ADD_11595

//ADD_8862 replaced by ADD_11602

//ADD_8861 replaced by ADD_11602

//BasicMUL48_165 replaced by BasicMUL48_970

//BasicMUL48_166 replaced by BasicMUL48_967

//BasicMUL48_167 replaced by BasicMUL48_970

//ADD_8866 replaced by ADD_11602

//ADD_8865 replaced by ADD_11602

//ADD_8864 replaced by ADD_11602

//ADD_8869 replaced by ADD_11601

//ADD_8868 replaced by ADD_11602

//ADD_8867 replaced by ADD_11602

//ADD_8871 replaced by ADD_11602

//ADD_8870 replaced by ADD_11602

//BasicMUL48_168 replaced by BasicMUL48_971

//BasicMUL48_169 replaced by BasicMUL48_970

//BasicMUL48_170 replaced by BasicMUL48_971

//ADD_8874 replaced by ADD_11595

//ADD_8873 replaced by ADD_11602

//ADD_8872 replaced by ADD_11602

//ADD_8877 replaced by ADD_11592

//ADD_8876 replaced by ADD_11602

//ADD_8875 replaced by ADD_11602

//ADD_8880 replaced by ADD_11592

//ADD_8879 replaced by ADD_11602

//ADD_8878 replaced by ADD_11602

//ADD_8883 replaced by ADD_11595

//ADD_8882 replaced by ADD_11602

//ADD_8881 replaced by ADD_11602

//BasicMUL48_171 replaced by BasicMUL48_970

//BasicMUL48_172 replaced by BasicMUL48_967

//BasicMUL48_173 replaced by BasicMUL48_970

//ADD_8886 replaced by ADD_11563

//ADD_8885 replaced by ADD_11602

//ADD_8884 replaced by ADD_11602

//ADD_8889 replaced by ADD_11560

//ADD_8888 replaced by ADD_11602

//ADD_8887 replaced by ADD_11602

//ADD_8892 replaced by ADD_11560

//ADD_8891 replaced by ADD_11602

//ADD_8890 replaced by ADD_11602

//ADD_8895 replaced by ADD_11563

//ADD_8894 replaced by ADD_11602

//ADD_8893 replaced by ADD_11602

//BasicMUL48_174 replaced by BasicMUL48_967

//BasicMUL48_175 replaced by BasicMUL48_958

//BasicMUL48_176 replaced by BasicMUL48_967

//ADD_8898 replaced by ADD_11595

//ADD_8897 replaced by ADD_11602

//ADD_8896 replaced by ADD_11602

//ADD_8901 replaced by ADD_11592

//ADD_8900 replaced by ADD_11602

//ADD_8899 replaced by ADD_11602

//ADD_8904 replaced by ADD_11592

//ADD_8903 replaced by ADD_11602

//ADD_8902 replaced by ADD_11602

//ADD_8907 replaced by ADD_11595

//ADD_8906 replaced by ADD_11602

//ADD_8905 replaced by ADD_11602

//BasicMUL48_177 replaced by BasicMUL48_970

//BasicMUL48_178 replaced by BasicMUL48_967

//BasicMUL48_179 replaced by BasicMUL48_970

//ADD_8910 replaced by ADD_11602

//ADD_8909 replaced by ADD_11602

//ADD_8908 replaced by ADD_11602

//ADD_8913 replaced by ADD_11601

//ADD_8912 replaced by ADD_11602

//ADD_8911 replaced by ADD_11602

//ADD_8915 replaced by ADD_11602

//ADD_8914 replaced by ADD_11602

//BasicMUL48_180 replaced by BasicMUL48_971

//BasicMUL48_181 replaced by BasicMUL48_970

//BasicMUL48_182 replaced by BasicMUL48_971

//ADD_8918 replaced by ADD_11595

//ADD_8917 replaced by ADD_11602

//ADD_8916 replaced by ADD_11602

//ADD_8921 replaced by ADD_11592

//ADD_8920 replaced by ADD_11602

//ADD_8919 replaced by ADD_11602

//ADD_8924 replaced by ADD_11592

//ADD_8923 replaced by ADD_11602

//ADD_8922 replaced by ADD_11602

//ADD_8927 replaced by ADD_11595

//ADD_8926 replaced by ADD_11602

//ADD_8925 replaced by ADD_11602

//BasicMUL48_183 replaced by BasicMUL48_970

//BasicMUL48_184 replaced by BasicMUL48_967

//BasicMUL48_185 replaced by BasicMUL48_970

//ADD_8930 replaced by ADD_11602

//ADD_8929 replaced by ADD_11602

//ADD_8928 replaced by ADD_11602

//ADD_8933 replaced by ADD_11601

//ADD_8932 replaced by ADD_11602

//ADD_8931 replaced by ADD_11602

//ADD_8935 replaced by ADD_11602

//ADD_8934 replaced by ADD_11602

//BasicMUL48_186 replaced by BasicMUL48_971

//BasicMUL48_187 replaced by BasicMUL48_970

//BasicMUL48_188 replaced by BasicMUL48_971

//ADD_8938 replaced by ADD_11602

//ADD_8937 replaced by ADD_11602

//ADD_8936 replaced by ADD_11602

//ADD_8941 replaced by ADD_11601

//ADD_8940 replaced by ADD_11602

//ADD_8939 replaced by ADD_11602

//ADD_8943 replaced by ADD_11602

//ADD_8942 replaced by ADD_11602

//BasicMUL48_189 replaced by BasicMUL48_971

//BasicMUL48_190 replaced by BasicMUL48_970

//BasicMUL48_191 replaced by BasicMUL48_971

//ADD_8946 replaced by ADD_11595

//ADD_8945 replaced by ADD_11602

//ADD_8944 replaced by ADD_11602

//ADD_8949 replaced by ADD_11592

//ADD_8948 replaced by ADD_11602

//ADD_8947 replaced by ADD_11602

//ADD_8952 replaced by ADD_11592

//ADD_8951 replaced by ADD_11602

//ADD_8950 replaced by ADD_11602

//ADD_8955 replaced by ADD_11595

//ADD_8954 replaced by ADD_11602

//ADD_8953 replaced by ADD_11602

//BasicMUL48_192 replaced by BasicMUL48_970

//BasicMUL48_193 replaced by BasicMUL48_967

//BasicMUL48_194 replaced by BasicMUL48_970

//ADD_8958 replaced by ADD_11602

//ADD_8957 replaced by ADD_11602

//ADD_8956 replaced by ADD_11602

//ADD_8961 replaced by ADD_11601

//ADD_8960 replaced by ADD_11602

//ADD_8959 replaced by ADD_11602

//ADD_8963 replaced by ADD_11602

//ADD_8962 replaced by ADD_11602

//BasicMUL48_195 replaced by BasicMUL48_971

//BasicMUL48_196 replaced by BasicMUL48_970

//BasicMUL48_197 replaced by BasicMUL48_971

//ADD_8966 replaced by ADD_11595

//ADD_8965 replaced by ADD_11602

//ADD_8964 replaced by ADD_11602

//ADD_8969 replaced by ADD_11592

//ADD_8968 replaced by ADD_11602

//ADD_8967 replaced by ADD_11602

//ADD_8972 replaced by ADD_11592

//ADD_8971 replaced by ADD_11602

//ADD_8970 replaced by ADD_11602

//ADD_8975 replaced by ADD_11595

//ADD_8974 replaced by ADD_11602

//ADD_8973 replaced by ADD_11602

//BasicMUL48_198 replaced by BasicMUL48_970

//BasicMUL48_199 replaced by BasicMUL48_967

//BasicMUL48_200 replaced by BasicMUL48_970

//ADD_8978 replaced by ADD_11563

//ADD_8977 replaced by ADD_11602

//ADD_8976 replaced by ADD_11602

//ADD_8981 replaced by ADD_11560

//ADD_8980 replaced by ADD_11602

//ADD_8979 replaced by ADD_11602

//ADD_8984 replaced by ADD_11560

//ADD_8983 replaced by ADD_11602

//ADD_8982 replaced by ADD_11602

//ADD_8987 replaced by ADD_11563

//ADD_8986 replaced by ADD_11602

//ADD_8985 replaced by ADD_11602

//BasicMUL48_201 replaced by BasicMUL48_967

//BasicMUL48_202 replaced by BasicMUL48_958

//BasicMUL48_203 replaced by BasicMUL48_967

//ADD_8990 replaced by ADD_11595

//ADD_8989 replaced by ADD_11602

//ADD_8988 replaced by ADD_11602

//ADD_8993 replaced by ADD_11592

//ADD_8992 replaced by ADD_11602

//ADD_8991 replaced by ADD_11602

//ADD_8996 replaced by ADD_11592

//ADD_8995 replaced by ADD_11602

//ADD_8994 replaced by ADD_11602

//ADD_8999 replaced by ADD_11595

//ADD_8998 replaced by ADD_11602

//ADD_8997 replaced by ADD_11602

//BasicMUL48_204 replaced by BasicMUL48_970

//BasicMUL48_205 replaced by BasicMUL48_967

//BasicMUL48_206 replaced by BasicMUL48_970

//ADD_9002 replaced by ADD_11602

//ADD_9001 replaced by ADD_11602

//ADD_9000 replaced by ADD_11602

//ADD_9005 replaced by ADD_11601

//ADD_9004 replaced by ADD_11602

//ADD_9003 replaced by ADD_11602

//ADD_9007 replaced by ADD_11602

//ADD_9006 replaced by ADD_11602

//BasicMUL48_207 replaced by BasicMUL48_971

//BasicMUL48_208 replaced by BasicMUL48_970

//BasicMUL48_209 replaced by BasicMUL48_971

//ADD_9010 replaced by ADD_11595

//ADD_9009 replaced by ADD_11602

//ADD_9008 replaced by ADD_11602

//ADD_9013 replaced by ADD_11592

//ADD_9012 replaced by ADD_11602

//ADD_9011 replaced by ADD_11602

//ADD_9016 replaced by ADD_11592

//ADD_9015 replaced by ADD_11602

//ADD_9014 replaced by ADD_11602

//ADD_9019 replaced by ADD_11595

//ADD_9018 replaced by ADD_11602

//ADD_9017 replaced by ADD_11602

//BasicMUL48_210 replaced by BasicMUL48_970

//BasicMUL48_211 replaced by BasicMUL48_967

//BasicMUL48_212 replaced by BasicMUL48_970

//ADD_9022 replaced by ADD_11602

//ADD_9021 replaced by ADD_11602

//ADD_9020 replaced by ADD_11602

//ADD_9025 replaced by ADD_11601

//ADD_9024 replaced by ADD_11602

//ADD_9023 replaced by ADD_11602

//ADD_9027 replaced by ADD_11602

//ADD_9026 replaced by ADD_11602

//BasicMUL48_213 replaced by BasicMUL48_971

//BasicMUL48_214 replaced by BasicMUL48_970

//BasicMUL48_215 replaced by BasicMUL48_971

//ADD_9030 replaced by ADD_11602

//ADD_9029 replaced by ADD_11602

//ADD_9028 replaced by ADD_11602

//ADD_9033 replaced by ADD_11601

//ADD_9032 replaced by ADD_11602

//ADD_9031 replaced by ADD_11602

//ADD_9035 replaced by ADD_11602

//ADD_9034 replaced by ADD_11602

//BasicMUL48_216 replaced by BasicMUL48_971

//BasicMUL48_217 replaced by BasicMUL48_970

//BasicMUL48_218 replaced by BasicMUL48_971

//ADD_9038 replaced by ADD_11595

//ADD_9037 replaced by ADD_11602

//ADD_9036 replaced by ADD_11602

//ADD_9041 replaced by ADD_11592

//ADD_9040 replaced by ADD_11602

//ADD_9039 replaced by ADD_11602

//ADD_9044 replaced by ADD_11592

//ADD_9043 replaced by ADD_11602

//ADD_9042 replaced by ADD_11602

//ADD_9047 replaced by ADD_11595

//ADD_9046 replaced by ADD_11602

//ADD_9045 replaced by ADD_11602

//BasicMUL48_219 replaced by BasicMUL48_970

//BasicMUL48_220 replaced by BasicMUL48_967

//BasicMUL48_221 replaced by BasicMUL48_970

//ADD_9050 replaced by ADD_11602

//ADD_9049 replaced by ADD_11602

//ADD_9048 replaced by ADD_11602

//ADD_9053 replaced by ADD_11601

//ADD_9052 replaced by ADD_11602

//ADD_9051 replaced by ADD_11602

//ADD_9055 replaced by ADD_11602

//ADD_9054 replaced by ADD_11602

//BasicMUL48_222 replaced by BasicMUL48_971

//BasicMUL48_223 replaced by BasicMUL48_970

//BasicMUL48_224 replaced by BasicMUL48_971

//ADD_9058 replaced by ADD_11595

//ADD_9057 replaced by ADD_11602

//ADD_9056 replaced by ADD_11602

//ADD_9061 replaced by ADD_11592

//ADD_9060 replaced by ADD_11602

//ADD_9059 replaced by ADD_11602

//ADD_9064 replaced by ADD_11592

//ADD_9063 replaced by ADD_11602

//ADD_9062 replaced by ADD_11602

//ADD_9067 replaced by ADD_11595

//ADD_9066 replaced by ADD_11602

//ADD_9065 replaced by ADD_11602

//BasicMUL48_225 replaced by BasicMUL48_970

//BasicMUL48_226 replaced by BasicMUL48_967

//BasicMUL48_227 replaced by BasicMUL48_970

//ADD_9070 replaced by ADD_11563

//ADD_9069 replaced by ADD_11602

//ADD_9068 replaced by ADD_11602

//ADD_9073 replaced by ADD_11560

//ADD_9072 replaced by ADD_11602

//ADD_9071 replaced by ADD_11602

//ADD_9076 replaced by ADD_11560

//ADD_9075 replaced by ADD_11602

//ADD_9074 replaced by ADD_11602

//ADD_9079 replaced by ADD_11563

//ADD_9078 replaced by ADD_11602

//ADD_9077 replaced by ADD_11602

//BasicMUL48_228 replaced by BasicMUL48_967

//BasicMUL48_229 replaced by BasicMUL48_958

//BasicMUL48_230 replaced by BasicMUL48_967

//ADD_9082 replaced by ADD_11595

//ADD_9081 replaced by ADD_11602

//ADD_9080 replaced by ADD_11602

//ADD_9085 replaced by ADD_11592

//ADD_9084 replaced by ADD_11602

//ADD_9083 replaced by ADD_11602

//ADD_9088 replaced by ADD_11592

//ADD_9087 replaced by ADD_11602

//ADD_9086 replaced by ADD_11602

//ADD_9091 replaced by ADD_11595

//ADD_9090 replaced by ADD_11602

//ADD_9089 replaced by ADD_11602

//BasicMUL48_231 replaced by BasicMUL48_970

//BasicMUL48_232 replaced by BasicMUL48_967

//BasicMUL48_233 replaced by BasicMUL48_970

//ADD_9094 replaced by ADD_11602

//ADD_9093 replaced by ADD_11602

//ADD_9092 replaced by ADD_11602

//ADD_9097 replaced by ADD_11601

//ADD_9096 replaced by ADD_11602

//ADD_9095 replaced by ADD_11602

//ADD_9099 replaced by ADD_11602

//ADD_9098 replaced by ADD_11602

//BasicMUL48_234 replaced by BasicMUL48_971

//BasicMUL48_235 replaced by BasicMUL48_970

//BasicMUL48_236 replaced by BasicMUL48_971

//ADD_9102 replaced by ADD_11595

//ADD_9101 replaced by ADD_11602

//ADD_9100 replaced by ADD_11602

//ADD_9105 replaced by ADD_11592

//ADD_9104 replaced by ADD_11602

//ADD_9103 replaced by ADD_11602

//ADD_9108 replaced by ADD_11592

//ADD_9107 replaced by ADD_11602

//ADD_9106 replaced by ADD_11602

//ADD_9111 replaced by ADD_11595

//ADD_9110 replaced by ADD_11602

//ADD_9109 replaced by ADD_11602

//BasicMUL48_237 replaced by BasicMUL48_970

//BasicMUL48_238 replaced by BasicMUL48_967

//BasicMUL48_239 replaced by BasicMUL48_970

//ADD_9114 replaced by ADD_11602

//ADD_9113 replaced by ADD_11602

//ADD_9112 replaced by ADD_11602

//ADD_9117 replaced by ADD_11601

//ADD_9116 replaced by ADD_11602

//ADD_9115 replaced by ADD_11602

//ADD_9119 replaced by ADD_11602

//ADD_9118 replaced by ADD_11602

//BasicMUL48_240 replaced by BasicMUL48_971

//BasicMUL48_241 replaced by BasicMUL48_970

//BasicMUL48_242 replaced by BasicMUL48_971

//ADD_9122 replaced by ADD_11602

//ADD_9121 replaced by ADD_11602

//ADD_9120 replaced by ADD_11602

//ADD_9125 replaced by ADD_11601

//ADD_9124 replaced by ADD_11602

//ADD_9123 replaced by ADD_11602

//ADD_9127 replaced by ADD_11602

//ADD_9126 replaced by ADD_11602

//BasicMUL48_243 replaced by BasicMUL48_971

//BasicMUL48_244 replaced by BasicMUL48_970

//BasicMUL48_245 replaced by BasicMUL48_971

//ADD_9130 replaced by ADD_11595

//ADD_9129 replaced by ADD_11602

//ADD_9128 replaced by ADD_11602

//ADD_9133 replaced by ADD_11592

//ADD_9132 replaced by ADD_11602

//ADD_9131 replaced by ADD_11602

//ADD_9136 replaced by ADD_11592

//ADD_9135 replaced by ADD_11602

//ADD_9134 replaced by ADD_11602

//ADD_9139 replaced by ADD_11595

//ADD_9138 replaced by ADD_11602

//ADD_9137 replaced by ADD_11602

//BasicMUL48_246 replaced by BasicMUL48_970

//BasicMUL48_247 replaced by BasicMUL48_967

//BasicMUL48_248 replaced by BasicMUL48_970

//ADD_9142 replaced by ADD_11602

//ADD_9141 replaced by ADD_11602

//ADD_9140 replaced by ADD_11602

//ADD_9145 replaced by ADD_11601

//ADD_9144 replaced by ADD_11602

//ADD_9143 replaced by ADD_11602

//ADD_9147 replaced by ADD_11602

//ADD_9146 replaced by ADD_11602

//BasicMUL48_249 replaced by BasicMUL48_971

//BasicMUL48_250 replaced by BasicMUL48_970

//BasicMUL48_251 replaced by BasicMUL48_971

//ADD_9150 replaced by ADD_11595

//ADD_9149 replaced by ADD_11602

//ADD_9148 replaced by ADD_11602

//ADD_9153 replaced by ADD_11592

//ADD_9152 replaced by ADD_11602

//ADD_9151 replaced by ADD_11602

//ADD_9156 replaced by ADD_11592

//ADD_9155 replaced by ADD_11602

//ADD_9154 replaced by ADD_11602

//ADD_9159 replaced by ADD_11595

//ADD_9158 replaced by ADD_11602

//ADD_9157 replaced by ADD_11602

//BasicMUL48_252 replaced by BasicMUL48_970

//BasicMUL48_253 replaced by BasicMUL48_967

//BasicMUL48_254 replaced by BasicMUL48_970

//ADD_9162 replaced by ADD_11563

//ADD_9161 replaced by ADD_11602

//ADD_9160 replaced by ADD_11602

//ADD_9165 replaced by ADD_11560

//ADD_9164 replaced by ADD_11602

//ADD_9163 replaced by ADD_11602

//ADD_9168 replaced by ADD_11560

//ADD_9167 replaced by ADD_11602

//ADD_9166 replaced by ADD_11602

//ADD_9171 replaced by ADD_11563

//ADD_9170 replaced by ADD_11602

//ADD_9169 replaced by ADD_11602

//BasicMUL48_255 replaced by BasicMUL48_967

//BasicMUL48_256 replaced by BasicMUL48_958

//BasicMUL48_257 replaced by BasicMUL48_967

//ADD_9174 replaced by ADD_11595

//ADD_9173 replaced by ADD_11602

//ADD_9172 replaced by ADD_11602

//ADD_9177 replaced by ADD_11592

//ADD_9176 replaced by ADD_11602

//ADD_9175 replaced by ADD_11602

//ADD_9180 replaced by ADD_11592

//ADD_9179 replaced by ADD_11602

//ADD_9178 replaced by ADD_11602

//ADD_9183 replaced by ADD_11595

//ADD_9182 replaced by ADD_11602

//ADD_9181 replaced by ADD_11602

//BasicMUL48_258 replaced by BasicMUL48_970

//BasicMUL48_259 replaced by BasicMUL48_967

//BasicMUL48_260 replaced by BasicMUL48_970

//ADD_9186 replaced by ADD_11602

//ADD_9185 replaced by ADD_11602

//ADD_9184 replaced by ADD_11602

//ADD_9189 replaced by ADD_11601

//ADD_9188 replaced by ADD_11602

//ADD_9187 replaced by ADD_11602

//ADD_9191 replaced by ADD_11602

//ADD_9190 replaced by ADD_11602

//BasicMUL48_261 replaced by BasicMUL48_971

//BasicMUL48_262 replaced by BasicMUL48_970

//BasicMUL48_263 replaced by BasicMUL48_971

//ADD_9194 replaced by ADD_11595

//ADD_9193 replaced by ADD_11602

//ADD_9192 replaced by ADD_11602

//ADD_9197 replaced by ADD_11592

//ADD_9196 replaced by ADD_11602

//ADD_9195 replaced by ADD_11602

//ADD_9200 replaced by ADD_11592

//ADD_9199 replaced by ADD_11602

//ADD_9198 replaced by ADD_11602

//ADD_9203 replaced by ADD_11595

//ADD_9202 replaced by ADD_11602

//ADD_9201 replaced by ADD_11602

//BasicMUL48_264 replaced by BasicMUL48_970

//BasicMUL48_265 replaced by BasicMUL48_967

//BasicMUL48_266 replaced by BasicMUL48_970

//ADD_9206 replaced by ADD_11602

//ADD_9205 replaced by ADD_11602

//ADD_9204 replaced by ADD_11602

//ADD_9209 replaced by ADD_11601

//ADD_9208 replaced by ADD_11602

//ADD_9207 replaced by ADD_11602

//ADD_9211 replaced by ADD_11602

//ADD_9210 replaced by ADD_11602

//BasicMUL48_267 replaced by BasicMUL48_971

//BasicMUL48_268 replaced by BasicMUL48_970

//BasicMUL48_269 replaced by BasicMUL48_971

//ADD_9214 replaced by ADD_11602

//ADD_9213 replaced by ADD_11602

//ADD_9212 replaced by ADD_11602

//ADD_9217 replaced by ADD_11601

//ADD_9216 replaced by ADD_11602

//ADD_9215 replaced by ADD_11602

//ADD_9219 replaced by ADD_11602

//ADD_9218 replaced by ADD_11602

//BasicMUL48_270 replaced by BasicMUL48_971

//BasicMUL48_271 replaced by BasicMUL48_970

//BasicMUL48_272 replaced by BasicMUL48_971

//ADD_9222 replaced by ADD_11595

//ADD_9221 replaced by ADD_11602

//ADD_9220 replaced by ADD_11602

//ADD_9225 replaced by ADD_11592

//ADD_9224 replaced by ADD_11602

//ADD_9223 replaced by ADD_11602

//ADD_9228 replaced by ADD_11592

//ADD_9227 replaced by ADD_11602

//ADD_9226 replaced by ADD_11602

//ADD_9231 replaced by ADD_11595

//ADD_9230 replaced by ADD_11602

//ADD_9229 replaced by ADD_11602

//BasicMUL48_273 replaced by BasicMUL48_970

//BasicMUL48_274 replaced by BasicMUL48_967

//BasicMUL48_275 replaced by BasicMUL48_970

//ADD_9234 replaced by ADD_11602

//ADD_9233 replaced by ADD_11602

//ADD_9232 replaced by ADD_11602

//ADD_9237 replaced by ADD_11601

//ADD_9236 replaced by ADD_11602

//ADD_9235 replaced by ADD_11602

//ADD_9239 replaced by ADD_11602

//ADD_9238 replaced by ADD_11602

//BasicMUL48_276 replaced by BasicMUL48_971

//BasicMUL48_277 replaced by BasicMUL48_970

//BasicMUL48_278 replaced by BasicMUL48_971

//ADD_9242 replaced by ADD_11595

//ADD_9241 replaced by ADD_11602

//ADD_9240 replaced by ADD_11602

//ADD_9245 replaced by ADD_11592

//ADD_9244 replaced by ADD_11602

//ADD_9243 replaced by ADD_11602

//ADD_9248 replaced by ADD_11592

//ADD_9247 replaced by ADD_11602

//ADD_9246 replaced by ADD_11602

//ADD_9251 replaced by ADD_11595

//ADD_9250 replaced by ADD_11602

//ADD_9249 replaced by ADD_11602

//BasicMUL48_279 replaced by BasicMUL48_970

//BasicMUL48_280 replaced by BasicMUL48_967

//BasicMUL48_281 replaced by BasicMUL48_970

//ADD_9254 replaced by ADD_11563

//ADD_9253 replaced by ADD_11602

//ADD_9252 replaced by ADD_11602

//ADD_9257 replaced by ADD_11560

//ADD_9256 replaced by ADD_11602

//ADD_9255 replaced by ADD_11602

//ADD_9260 replaced by ADD_11560

//ADD_9259 replaced by ADD_11602

//ADD_9258 replaced by ADD_11602

//ADD_9263 replaced by ADD_11563

//ADD_9262 replaced by ADD_11602

//ADD_9261 replaced by ADD_11602

//BasicMUL48_282 replaced by BasicMUL48_967

//BasicMUL48_283 replaced by BasicMUL48_958

//BasicMUL48_284 replaced by BasicMUL48_967

//ADD_9266 replaced by ADD_11595

//ADD_9265 replaced by ADD_11602

//ADD_9264 replaced by ADD_11602

//ADD_9269 replaced by ADD_11592

//ADD_9268 replaced by ADD_11602

//ADD_9267 replaced by ADD_11602

//ADD_9272 replaced by ADD_11592

//ADD_9271 replaced by ADD_11602

//ADD_9270 replaced by ADD_11602

//ADD_9275 replaced by ADD_11595

//ADD_9274 replaced by ADD_11602

//ADD_9273 replaced by ADD_11602

//BasicMUL48_285 replaced by BasicMUL48_970

//BasicMUL48_286 replaced by BasicMUL48_967

//BasicMUL48_287 replaced by BasicMUL48_970

//ADD_9278 replaced by ADD_11602

//ADD_9277 replaced by ADD_11602

//ADD_9276 replaced by ADD_11602

//ADD_9281 replaced by ADD_11601

//ADD_9280 replaced by ADD_11602

//ADD_9279 replaced by ADD_11602

//ADD_9283 replaced by ADD_11602

//ADD_9282 replaced by ADD_11602

//BasicMUL48_288 replaced by BasicMUL48_971

//BasicMUL48_289 replaced by BasicMUL48_970

//BasicMUL48_290 replaced by BasicMUL48_971

//ADD_9286 replaced by ADD_11595

//ADD_9285 replaced by ADD_11602

//ADD_9284 replaced by ADD_11602

//ADD_9289 replaced by ADD_11592

//ADD_9288 replaced by ADD_11602

//ADD_9287 replaced by ADD_11602

//ADD_9292 replaced by ADD_11592

//ADD_9291 replaced by ADD_11602

//ADD_9290 replaced by ADD_11602

//ADD_9295 replaced by ADD_11595

//ADD_9294 replaced by ADD_11602

//ADD_9293 replaced by ADD_11602

//BasicMUL48_291 replaced by BasicMUL48_970

//BasicMUL48_292 replaced by BasicMUL48_967

//BasicMUL48_293 replaced by BasicMUL48_970

//ADD_9298 replaced by ADD_11602

//ADD_9297 replaced by ADD_11602

//ADD_9296 replaced by ADD_11602

//ADD_9301 replaced by ADD_11601

//ADD_9300 replaced by ADD_11602

//ADD_9299 replaced by ADD_11602

//ADD_9303 replaced by ADD_11602

//ADD_9302 replaced by ADD_11602

//BasicMUL48_294 replaced by BasicMUL48_971

//BasicMUL48_295 replaced by BasicMUL48_970

//BasicMUL48_296 replaced by BasicMUL48_971

//ADD_9306 replaced by ADD_11602

//ADD_9305 replaced by ADD_11602

//ADD_9304 replaced by ADD_11602

//ADD_9309 replaced by ADD_11601

//ADD_9308 replaced by ADD_11602

//ADD_9307 replaced by ADD_11602

//ADD_9311 replaced by ADD_11602

//ADD_9310 replaced by ADD_11602

//BasicMUL48_297 replaced by BasicMUL48_971

//BasicMUL48_298 replaced by BasicMUL48_970

//BasicMUL48_299 replaced by BasicMUL48_971

//ADD_9314 replaced by ADD_11595

//ADD_9313 replaced by ADD_11602

//ADD_9312 replaced by ADD_11602

//ADD_9317 replaced by ADD_11592

//ADD_9316 replaced by ADD_11602

//ADD_9315 replaced by ADD_11602

//ADD_9320 replaced by ADD_11592

//ADD_9319 replaced by ADD_11602

//ADD_9318 replaced by ADD_11602

//ADD_9323 replaced by ADD_11595

//ADD_9322 replaced by ADD_11602

//ADD_9321 replaced by ADD_11602

//BasicMUL48_300 replaced by BasicMUL48_970

//BasicMUL48_301 replaced by BasicMUL48_967

//BasicMUL48_302 replaced by BasicMUL48_970

//ADD_9326 replaced by ADD_11602

//ADD_9325 replaced by ADD_11602

//ADD_9324 replaced by ADD_11602

//ADD_9329 replaced by ADD_11601

//ADD_9328 replaced by ADD_11602

//ADD_9327 replaced by ADD_11602

//ADD_9331 replaced by ADD_11602

//ADD_9330 replaced by ADD_11602

//BasicMUL48_303 replaced by BasicMUL48_971

//BasicMUL48_304 replaced by BasicMUL48_970

//BasicMUL48_305 replaced by BasicMUL48_971

//ADD_9334 replaced by ADD_11595

//ADD_9333 replaced by ADD_11602

//ADD_9332 replaced by ADD_11602

//ADD_9337 replaced by ADD_11592

//ADD_9336 replaced by ADD_11602

//ADD_9335 replaced by ADD_11602

//ADD_9340 replaced by ADD_11592

//ADD_9339 replaced by ADD_11602

//ADD_9338 replaced by ADD_11602

//ADD_9343 replaced by ADD_11595

//ADD_9342 replaced by ADD_11602

//ADD_9341 replaced by ADD_11602

//BasicMUL48_306 replaced by BasicMUL48_970

//BasicMUL48_307 replaced by BasicMUL48_967

//BasicMUL48_308 replaced by BasicMUL48_970

//ADD_9346 replaced by ADD_11563

//ADD_9345 replaced by ADD_11602

//ADD_9344 replaced by ADD_11602

//ADD_9349 replaced by ADD_11560

//ADD_9348 replaced by ADD_11602

//ADD_9347 replaced by ADD_11602

//ADD_9352 replaced by ADD_11560

//ADD_9351 replaced by ADD_11602

//ADD_9350 replaced by ADD_11602

//ADD_9355 replaced by ADD_11563

//ADD_9354 replaced by ADD_11602

//ADD_9353 replaced by ADD_11602

//BasicMUL48_309 replaced by BasicMUL48_967

//BasicMUL48_310 replaced by BasicMUL48_958

//BasicMUL48_311 replaced by BasicMUL48_967

//ADD_9358 replaced by ADD_11595

//ADD_9357 replaced by ADD_11602

//ADD_9356 replaced by ADD_11602

//ADD_9361 replaced by ADD_11592

//ADD_9360 replaced by ADD_11602

//ADD_9359 replaced by ADD_11602

//ADD_9364 replaced by ADD_11592

//ADD_9363 replaced by ADD_11602

//ADD_9362 replaced by ADD_11602

//ADD_9367 replaced by ADD_11595

//ADD_9366 replaced by ADD_11602

//ADD_9365 replaced by ADD_11602

//BasicMUL48_312 replaced by BasicMUL48_970

//BasicMUL48_313 replaced by BasicMUL48_967

//BasicMUL48_314 replaced by BasicMUL48_970

//ADD_9370 replaced by ADD_11602

//ADD_9369 replaced by ADD_11602

//ADD_9368 replaced by ADD_11602

//ADD_9373 replaced by ADD_11601

//ADD_9372 replaced by ADD_11602

//ADD_9371 replaced by ADD_11602

//ADD_9375 replaced by ADD_11602

//ADD_9374 replaced by ADD_11602

//BasicMUL48_315 replaced by BasicMUL48_971

//BasicMUL48_316 replaced by BasicMUL48_970

//BasicMUL48_317 replaced by BasicMUL48_971

//ADD_9378 replaced by ADD_11595

//ADD_9377 replaced by ADD_11602

//ADD_9376 replaced by ADD_11602

//ADD_9381 replaced by ADD_11592

//ADD_9380 replaced by ADD_11602

//ADD_9379 replaced by ADD_11602

//ADD_9384 replaced by ADD_11592

//ADD_9383 replaced by ADD_11602

//ADD_9382 replaced by ADD_11602

//ADD_9387 replaced by ADD_11595

//ADD_9386 replaced by ADD_11602

//ADD_9385 replaced by ADD_11602

//BasicMUL48_318 replaced by BasicMUL48_970

//BasicMUL48_319 replaced by BasicMUL48_967

//BasicMUL48_320 replaced by BasicMUL48_970

//ADD_9390 replaced by ADD_11602

//ADD_9389 replaced by ADD_11602

//ADD_9388 replaced by ADD_11602

//ADD_9393 replaced by ADD_11601

//ADD_9392 replaced by ADD_11602

//ADD_9391 replaced by ADD_11602

//ADD_9395 replaced by ADD_11602

//ADD_9394 replaced by ADD_11602

//BasicMUL48_321 replaced by BasicMUL48_971

//BasicMUL48_322 replaced by BasicMUL48_970

//BasicMUL48_323 replaced by BasicMUL48_971

//ADD_9398 replaced by ADD_11602

//ADD_9397 replaced by ADD_11602

//ADD_9396 replaced by ADD_11602

//ADD_9401 replaced by ADD_11601

//ADD_9400 replaced by ADD_11602

//ADD_9399 replaced by ADD_11602

//ADD_9403 replaced by ADD_11602

//ADD_9402 replaced by ADD_11602

//BasicMUL48_324 replaced by BasicMUL48_971

//BasicMUL48_325 replaced by BasicMUL48_970

//BasicMUL48_326 replaced by BasicMUL48_971

//ADD_9406 replaced by ADD_11595

//ADD_9405 replaced by ADD_11602

//ADD_9404 replaced by ADD_11602

//ADD_9409 replaced by ADD_11592

//ADD_9408 replaced by ADD_11602

//ADD_9407 replaced by ADD_11602

//ADD_9412 replaced by ADD_11592

//ADD_9411 replaced by ADD_11602

//ADD_9410 replaced by ADD_11602

//ADD_9415 replaced by ADD_11595

//ADD_9414 replaced by ADD_11602

//ADD_9413 replaced by ADD_11602

//BasicMUL48_327 replaced by BasicMUL48_970

//BasicMUL48_328 replaced by BasicMUL48_967

//BasicMUL48_329 replaced by BasicMUL48_970

//ADD_9418 replaced by ADD_11602

//ADD_9417 replaced by ADD_11602

//ADD_9416 replaced by ADD_11602

//ADD_9421 replaced by ADD_11601

//ADD_9420 replaced by ADD_11602

//ADD_9419 replaced by ADD_11602

//ADD_9423 replaced by ADD_11602

//ADD_9422 replaced by ADD_11602

//BasicMUL48_330 replaced by BasicMUL48_971

//BasicMUL48_331 replaced by BasicMUL48_970

//BasicMUL48_332 replaced by BasicMUL48_971

//ADD_9426 replaced by ADD_11595

//ADD_9425 replaced by ADD_11602

//ADD_9424 replaced by ADD_11602

//ADD_9429 replaced by ADD_11592

//ADD_9428 replaced by ADD_11602

//ADD_9427 replaced by ADD_11602

//ADD_9432 replaced by ADD_11592

//ADD_9431 replaced by ADD_11602

//ADD_9430 replaced by ADD_11602

//ADD_9435 replaced by ADD_11595

//ADD_9434 replaced by ADD_11602

//ADD_9433 replaced by ADD_11602

//BasicMUL48_333 replaced by BasicMUL48_970

//BasicMUL48_334 replaced by BasicMUL48_967

//BasicMUL48_335 replaced by BasicMUL48_970

//ADD_9438 replaced by ADD_11563

//ADD_9437 replaced by ADD_11602

//ADD_9436 replaced by ADD_11602

//ADD_9441 replaced by ADD_11560

//ADD_9440 replaced by ADD_11602

//ADD_9439 replaced by ADD_11602

//ADD_9444 replaced by ADD_11560

//ADD_9443 replaced by ADD_11602

//ADD_9442 replaced by ADD_11602

//ADD_9447 replaced by ADD_11563

//ADD_9446 replaced by ADD_11602

//ADD_9445 replaced by ADD_11602

//BasicMUL48_336 replaced by BasicMUL48_967

//BasicMUL48_337 replaced by BasicMUL48_958

//BasicMUL48_338 replaced by BasicMUL48_967

//ADD_9450 replaced by ADD_11595

//ADD_9449 replaced by ADD_11602

//ADD_9448 replaced by ADD_11602

//ADD_9453 replaced by ADD_11592

//ADD_9452 replaced by ADD_11602

//ADD_9451 replaced by ADD_11602

//ADD_9456 replaced by ADD_11592

//ADD_9455 replaced by ADD_11602

//ADD_9454 replaced by ADD_11602

//ADD_9459 replaced by ADD_11595

//ADD_9458 replaced by ADD_11602

//ADD_9457 replaced by ADD_11602

//BasicMUL48_339 replaced by BasicMUL48_970

//BasicMUL48_340 replaced by BasicMUL48_967

//BasicMUL48_341 replaced by BasicMUL48_970

//ADD_9462 replaced by ADD_11602

//ADD_9461 replaced by ADD_11602

//ADD_9460 replaced by ADD_11602

//ADD_9465 replaced by ADD_11601

//ADD_9464 replaced by ADD_11602

//ADD_9463 replaced by ADD_11602

//ADD_9467 replaced by ADD_11602

//ADD_9466 replaced by ADD_11602

//BasicMUL48_342 replaced by BasicMUL48_971

//BasicMUL48_343 replaced by BasicMUL48_970

//BasicMUL48_344 replaced by BasicMUL48_971

//ADD_9470 replaced by ADD_11595

//ADD_9469 replaced by ADD_11602

//ADD_9468 replaced by ADD_11602

//ADD_9473 replaced by ADD_11592

//ADD_9472 replaced by ADD_11602

//ADD_9471 replaced by ADD_11602

//ADD_9476 replaced by ADD_11592

//ADD_9475 replaced by ADD_11602

//ADD_9474 replaced by ADD_11602

//ADD_9479 replaced by ADD_11595

//ADD_9478 replaced by ADD_11602

//ADD_9477 replaced by ADD_11602

//BasicMUL48_345 replaced by BasicMUL48_970

//BasicMUL48_346 replaced by BasicMUL48_967

//BasicMUL48_347 replaced by BasicMUL48_970

//ADD_9482 replaced by ADD_11602

//ADD_9481 replaced by ADD_11602

//ADD_9480 replaced by ADD_11602

//ADD_9485 replaced by ADD_11601

//ADD_9484 replaced by ADD_11602

//ADD_9483 replaced by ADD_11602

//ADD_9487 replaced by ADD_11602

//ADD_9486 replaced by ADD_11602

//BasicMUL48_348 replaced by BasicMUL48_971

//BasicMUL48_349 replaced by BasicMUL48_970

//BasicMUL48_350 replaced by BasicMUL48_971

//ADD_9490 replaced by ADD_11602

//ADD_9489 replaced by ADD_11602

//ADD_9488 replaced by ADD_11602

//ADD_9493 replaced by ADD_11601

//ADD_9492 replaced by ADD_11602

//ADD_9491 replaced by ADD_11602

//ADD_9495 replaced by ADD_11602

//ADD_9494 replaced by ADD_11602

//BasicMUL48_351 replaced by BasicMUL48_971

//BasicMUL48_352 replaced by BasicMUL48_970

//BasicMUL48_353 replaced by BasicMUL48_971

//ADD_9498 replaced by ADD_11595

//ADD_9497 replaced by ADD_11602

//ADD_9496 replaced by ADD_11602

//ADD_9501 replaced by ADD_11592

//ADD_9500 replaced by ADD_11602

//ADD_9499 replaced by ADD_11602

//ADD_9504 replaced by ADD_11592

//ADD_9503 replaced by ADD_11602

//ADD_9502 replaced by ADD_11602

//ADD_9507 replaced by ADD_11595

//ADD_9506 replaced by ADD_11602

//ADD_9505 replaced by ADD_11602

//BasicMUL48_354 replaced by BasicMUL48_970

//BasicMUL48_355 replaced by BasicMUL48_967

//BasicMUL48_356 replaced by BasicMUL48_970

//ADD_9510 replaced by ADD_11602

//ADD_9509 replaced by ADD_11602

//ADD_9508 replaced by ADD_11602

//ADD_9513 replaced by ADD_11601

//ADD_9512 replaced by ADD_11602

//ADD_9511 replaced by ADD_11602

//ADD_9515 replaced by ADD_11602

//ADD_9514 replaced by ADD_11602

//BasicMUL48_357 replaced by BasicMUL48_971

//BasicMUL48_358 replaced by BasicMUL48_970

//BasicMUL48_359 replaced by BasicMUL48_971

//ADD_9518 replaced by ADD_11595

//ADD_9517 replaced by ADD_11602

//ADD_9516 replaced by ADD_11602

//ADD_9521 replaced by ADD_11592

//ADD_9520 replaced by ADD_11602

//ADD_9519 replaced by ADD_11602

//ADD_9524 replaced by ADD_11592

//ADD_9523 replaced by ADD_11602

//ADD_9522 replaced by ADD_11602

//ADD_9527 replaced by ADD_11595

//ADD_9526 replaced by ADD_11602

//ADD_9525 replaced by ADD_11602

//BasicMUL48_360 replaced by BasicMUL48_970

//BasicMUL48_361 replaced by BasicMUL48_967

//BasicMUL48_362 replaced by BasicMUL48_970

//ADD_9530 replaced by ADD_11563

//ADD_9529 replaced by ADD_11602

//ADD_9528 replaced by ADD_11602

//ADD_9533 replaced by ADD_11560

//ADD_9532 replaced by ADD_11602

//ADD_9531 replaced by ADD_11602

//ADD_9536 replaced by ADD_11560

//ADD_9535 replaced by ADD_11602

//ADD_9534 replaced by ADD_11602

//ADD_9539 replaced by ADD_11563

//ADD_9538 replaced by ADD_11602

//ADD_9537 replaced by ADD_11602

//BasicMUL48_363 replaced by BasicMUL48_967

//BasicMUL48_364 replaced by BasicMUL48_958

//BasicMUL48_365 replaced by BasicMUL48_967

//ADD_9542 replaced by ADD_11595

//ADD_9541 replaced by ADD_11602

//ADD_9540 replaced by ADD_11602

//ADD_9545 replaced by ADD_11592

//ADD_9544 replaced by ADD_11602

//ADD_9543 replaced by ADD_11602

//ADD_9548 replaced by ADD_11592

//ADD_9547 replaced by ADD_11602

//ADD_9546 replaced by ADD_11602

//ADD_9551 replaced by ADD_11595

//ADD_9550 replaced by ADD_11602

//ADD_9549 replaced by ADD_11602

//BasicMUL48_366 replaced by BasicMUL48_970

//BasicMUL48_367 replaced by BasicMUL48_967

//BasicMUL48_368 replaced by BasicMUL48_970

//ADD_9554 replaced by ADD_11602

//ADD_9553 replaced by ADD_11602

//ADD_9552 replaced by ADD_11602

//ADD_9557 replaced by ADD_11601

//ADD_9556 replaced by ADD_11602

//ADD_9555 replaced by ADD_11602

//ADD_9559 replaced by ADD_11602

//ADD_9558 replaced by ADD_11602

//BasicMUL48_369 replaced by BasicMUL48_971

//BasicMUL48_370 replaced by BasicMUL48_970

//BasicMUL48_371 replaced by BasicMUL48_971

//ADD_9562 replaced by ADD_11595

//ADD_9561 replaced by ADD_11602

//ADD_9560 replaced by ADD_11602

//ADD_9565 replaced by ADD_11592

//ADD_9564 replaced by ADD_11602

//ADD_9563 replaced by ADD_11602

//ADD_9568 replaced by ADD_11592

//ADD_9567 replaced by ADD_11602

//ADD_9566 replaced by ADD_11602

//ADD_9571 replaced by ADD_11595

//ADD_9570 replaced by ADD_11602

//ADD_9569 replaced by ADD_11602

//BasicMUL48_372 replaced by BasicMUL48_970

//BasicMUL48_373 replaced by BasicMUL48_967

//BasicMUL48_374 replaced by BasicMUL48_970

//ADD_9574 replaced by ADD_11602

//ADD_9573 replaced by ADD_11602

//ADD_9572 replaced by ADD_11602

//ADD_9577 replaced by ADD_11601

//ADD_9576 replaced by ADD_11602

//ADD_9575 replaced by ADD_11602

//ADD_9579 replaced by ADD_11602

//ADD_9578 replaced by ADD_11602

//BasicMUL48_375 replaced by BasicMUL48_971

//BasicMUL48_376 replaced by BasicMUL48_970

//BasicMUL48_377 replaced by BasicMUL48_971

//ADD_9582 replaced by ADD_11602

//ADD_9581 replaced by ADD_11602

//ADD_9580 replaced by ADD_11602

//ADD_9585 replaced by ADD_11601

//ADD_9584 replaced by ADD_11602

//ADD_9583 replaced by ADD_11602

//ADD_9587 replaced by ADD_11602

//ADD_9586 replaced by ADD_11602

//BasicMUL48_378 replaced by BasicMUL48_971

//BasicMUL48_379 replaced by BasicMUL48_970

//BasicMUL48_380 replaced by BasicMUL48_971

//ADD_9590 replaced by ADD_11595

//ADD_9589 replaced by ADD_11602

//ADD_9588 replaced by ADD_11602

//ADD_9593 replaced by ADD_11592

//ADD_9592 replaced by ADD_11602

//ADD_9591 replaced by ADD_11602

//ADD_9596 replaced by ADD_11592

//ADD_9595 replaced by ADD_11602

//ADD_9594 replaced by ADD_11602

//ADD_9599 replaced by ADD_11595

//ADD_9598 replaced by ADD_11602

//ADD_9597 replaced by ADD_11602

//BasicMUL48_381 replaced by BasicMUL48_970

//BasicMUL48_382 replaced by BasicMUL48_967

//BasicMUL48_383 replaced by BasicMUL48_970

//ADD_9602 replaced by ADD_11602

//ADD_9601 replaced by ADD_11602

//ADD_9600 replaced by ADD_11602

//ADD_9605 replaced by ADD_11601

//ADD_9604 replaced by ADD_11602

//ADD_9603 replaced by ADD_11602

//ADD_9607 replaced by ADD_11602

//ADD_9606 replaced by ADD_11602

//BasicMUL48_384 replaced by BasicMUL48_971

//BasicMUL48_385 replaced by BasicMUL48_970

//BasicMUL48_386 replaced by BasicMUL48_971

//ADD_9610 replaced by ADD_11595

//ADD_9609 replaced by ADD_11602

//ADD_9608 replaced by ADD_11602

//ADD_9613 replaced by ADD_11592

//ADD_9612 replaced by ADD_11602

//ADD_9611 replaced by ADD_11602

//ADD_9616 replaced by ADD_11592

//ADD_9615 replaced by ADD_11602

//ADD_9614 replaced by ADD_11602

//ADD_9619 replaced by ADD_11595

//ADD_9618 replaced by ADD_11602

//ADD_9617 replaced by ADD_11602

//BasicMUL48_387 replaced by BasicMUL48_970

//BasicMUL48_388 replaced by BasicMUL48_967

//BasicMUL48_389 replaced by BasicMUL48_970

//ADD_9622 replaced by ADD_11563

//ADD_9621 replaced by ADD_11602

//ADD_9620 replaced by ADD_11602

//ADD_9625 replaced by ADD_11560

//ADD_9624 replaced by ADD_11602

//ADD_9623 replaced by ADD_11602

//ADD_9628 replaced by ADD_11560

//ADD_9627 replaced by ADD_11602

//ADD_9626 replaced by ADD_11602

//ADD_9631 replaced by ADD_11563

//ADD_9630 replaced by ADD_11602

//ADD_9629 replaced by ADD_11602

//BasicMUL48_390 replaced by BasicMUL48_967

//BasicMUL48_391 replaced by BasicMUL48_958

//BasicMUL48_392 replaced by BasicMUL48_967

//ADD_9634 replaced by ADD_11595

//ADD_9633 replaced by ADD_11602

//ADD_9632 replaced by ADD_11602

//ADD_9637 replaced by ADD_11592

//ADD_9636 replaced by ADD_11602

//ADD_9635 replaced by ADD_11602

//ADD_9640 replaced by ADD_11592

//ADD_9639 replaced by ADD_11602

//ADD_9638 replaced by ADD_11602

//ADD_9643 replaced by ADD_11595

//ADD_9642 replaced by ADD_11602

//ADD_9641 replaced by ADD_11602

//BasicMUL48_393 replaced by BasicMUL48_970

//BasicMUL48_394 replaced by BasicMUL48_967

//BasicMUL48_395 replaced by BasicMUL48_970

//ADD_9646 replaced by ADD_11602

//ADD_9645 replaced by ADD_11602

//ADD_9644 replaced by ADD_11602

//ADD_9649 replaced by ADD_11601

//ADD_9648 replaced by ADD_11602

//ADD_9647 replaced by ADD_11602

//ADD_9651 replaced by ADD_11602

//ADD_9650 replaced by ADD_11602

//BasicMUL48_396 replaced by BasicMUL48_971

//BasicMUL48_397 replaced by BasicMUL48_970

//BasicMUL48_398 replaced by BasicMUL48_971

//ADD_9654 replaced by ADD_11595

//ADD_9653 replaced by ADD_11602

//ADD_9652 replaced by ADD_11602

//ADD_9657 replaced by ADD_11592

//ADD_9656 replaced by ADD_11602

//ADD_9655 replaced by ADD_11602

//ADD_9660 replaced by ADD_11592

//ADD_9659 replaced by ADD_11602

//ADD_9658 replaced by ADD_11602

//ADD_9663 replaced by ADD_11595

//ADD_9662 replaced by ADD_11602

//ADD_9661 replaced by ADD_11602

//BasicMUL48_399 replaced by BasicMUL48_970

//BasicMUL48_400 replaced by BasicMUL48_967

//BasicMUL48_401 replaced by BasicMUL48_970

//ADD_9666 replaced by ADD_11602

//ADD_9665 replaced by ADD_11602

//ADD_9664 replaced by ADD_11602

//ADD_9669 replaced by ADD_11601

//ADD_9668 replaced by ADD_11602

//ADD_9667 replaced by ADD_11602

//ADD_9671 replaced by ADD_11602

//ADD_9670 replaced by ADD_11602

//BasicMUL48_402 replaced by BasicMUL48_971

//BasicMUL48_403 replaced by BasicMUL48_970

//BasicMUL48_404 replaced by BasicMUL48_971

//ADD_9674 replaced by ADD_11602

//ADD_9673 replaced by ADD_11602

//ADD_9672 replaced by ADD_11602

//ADD_9677 replaced by ADD_11601

//ADD_9676 replaced by ADD_11602

//ADD_9675 replaced by ADD_11602

//ADD_9679 replaced by ADD_11602

//ADD_9678 replaced by ADD_11602

//BasicMUL48_405 replaced by BasicMUL48_971

//BasicMUL48_406 replaced by BasicMUL48_970

//BasicMUL48_407 replaced by BasicMUL48_971

//ADD_9682 replaced by ADD_11595

//ADD_9681 replaced by ADD_11602

//ADD_9680 replaced by ADD_11602

//ADD_9685 replaced by ADD_11592

//ADD_9684 replaced by ADD_11602

//ADD_9683 replaced by ADD_11602

//ADD_9688 replaced by ADD_11592

//ADD_9687 replaced by ADD_11602

//ADD_9686 replaced by ADD_11602

//ADD_9691 replaced by ADD_11595

//ADD_9690 replaced by ADD_11602

//ADD_9689 replaced by ADD_11602

//BasicMUL48_408 replaced by BasicMUL48_970

//BasicMUL48_409 replaced by BasicMUL48_967

//BasicMUL48_410 replaced by BasicMUL48_970

//ADD_9694 replaced by ADD_11602

//ADD_9693 replaced by ADD_11602

//ADD_9692 replaced by ADD_11602

//ADD_9697 replaced by ADD_11601

//ADD_9696 replaced by ADD_11602

//ADD_9695 replaced by ADD_11602

//ADD_9699 replaced by ADD_11602

//ADD_9698 replaced by ADD_11602

//BasicMUL48_411 replaced by BasicMUL48_971

//BasicMUL48_412 replaced by BasicMUL48_970

//BasicMUL48_413 replaced by BasicMUL48_971

//ADD_9702 replaced by ADD_11595

//ADD_9701 replaced by ADD_11602

//ADD_9700 replaced by ADD_11602

//ADD_9705 replaced by ADD_11592

//ADD_9704 replaced by ADD_11602

//ADD_9703 replaced by ADD_11602

//ADD_9708 replaced by ADD_11592

//ADD_9707 replaced by ADD_11602

//ADD_9706 replaced by ADD_11602

//ADD_9711 replaced by ADD_11595

//ADD_9710 replaced by ADD_11602

//ADD_9709 replaced by ADD_11602

//BasicMUL48_414 replaced by BasicMUL48_970

//BasicMUL48_415 replaced by BasicMUL48_967

//BasicMUL48_416 replaced by BasicMUL48_970

//ADD_9714 replaced by ADD_11563

//ADD_9713 replaced by ADD_11602

//ADD_9712 replaced by ADD_11602

//ADD_9717 replaced by ADD_11560

//ADD_9716 replaced by ADD_11602

//ADD_9715 replaced by ADD_11602

//ADD_9720 replaced by ADD_11560

//ADD_9719 replaced by ADD_11602

//ADD_9718 replaced by ADD_11602

//ADD_9723 replaced by ADD_11563

//ADD_9722 replaced by ADD_11602

//ADD_9721 replaced by ADD_11602

//BasicMUL48_417 replaced by BasicMUL48_967

//BasicMUL48_418 replaced by BasicMUL48_958

//BasicMUL48_419 replaced by BasicMUL48_967

//ADD_9726 replaced by ADD_11595

//ADD_9725 replaced by ADD_11602

//ADD_9724 replaced by ADD_11602

//ADD_9729 replaced by ADD_11592

//ADD_9728 replaced by ADD_11602

//ADD_9727 replaced by ADD_11602

//ADD_9732 replaced by ADD_11592

//ADD_9731 replaced by ADD_11602

//ADD_9730 replaced by ADD_11602

//ADD_9735 replaced by ADD_11595

//ADD_9734 replaced by ADD_11602

//ADD_9733 replaced by ADD_11602

//BasicMUL48_420 replaced by BasicMUL48_970

//BasicMUL48_421 replaced by BasicMUL48_967

//BasicMUL48_422 replaced by BasicMUL48_970

//ADD_9738 replaced by ADD_11602

//ADD_9737 replaced by ADD_11602

//ADD_9736 replaced by ADD_11602

//ADD_9741 replaced by ADD_11601

//ADD_9740 replaced by ADD_11602

//ADD_9739 replaced by ADD_11602

//ADD_9743 replaced by ADD_11602

//ADD_9742 replaced by ADD_11602

//BasicMUL48_423 replaced by BasicMUL48_971

//BasicMUL48_424 replaced by BasicMUL48_970

//BasicMUL48_425 replaced by BasicMUL48_971

//ADD_9746 replaced by ADD_11595

//ADD_9745 replaced by ADD_11602

//ADD_9744 replaced by ADD_11602

//ADD_9749 replaced by ADD_11592

//ADD_9748 replaced by ADD_11602

//ADD_9747 replaced by ADD_11602

//ADD_9752 replaced by ADD_11592

//ADD_9751 replaced by ADD_11602

//ADD_9750 replaced by ADD_11602

//ADD_9755 replaced by ADD_11595

//ADD_9754 replaced by ADD_11602

//ADD_9753 replaced by ADD_11602

//BasicMUL48_426 replaced by BasicMUL48_970

//BasicMUL48_427 replaced by BasicMUL48_967

//BasicMUL48_428 replaced by BasicMUL48_970

//ADD_9758 replaced by ADD_11602

//ADD_9757 replaced by ADD_11602

//ADD_9756 replaced by ADD_11602

//ADD_9761 replaced by ADD_11601

//ADD_9760 replaced by ADD_11602

//ADD_9759 replaced by ADD_11602

//ADD_9763 replaced by ADD_11602

//ADD_9762 replaced by ADD_11602

//BasicMUL48_429 replaced by BasicMUL48_971

//BasicMUL48_430 replaced by BasicMUL48_970

//BasicMUL48_431 replaced by BasicMUL48_971

//ADD_9766 replaced by ADD_11602

//ADD_9765 replaced by ADD_11602

//ADD_9764 replaced by ADD_11602

//ADD_9769 replaced by ADD_11601

//ADD_9768 replaced by ADD_11602

//ADD_9767 replaced by ADD_11602

//ADD_9771 replaced by ADD_11602

//ADD_9770 replaced by ADD_11602

//BasicMUL48_432 replaced by BasicMUL48_971

//BasicMUL48_433 replaced by BasicMUL48_970

//BasicMUL48_434 replaced by BasicMUL48_971

//ADD_9774 replaced by ADD_11595

//ADD_9773 replaced by ADD_11602

//ADD_9772 replaced by ADD_11602

//ADD_9777 replaced by ADD_11592

//ADD_9776 replaced by ADD_11602

//ADD_9775 replaced by ADD_11602

//ADD_9780 replaced by ADD_11592

//ADD_9779 replaced by ADD_11602

//ADD_9778 replaced by ADD_11602

//ADD_9783 replaced by ADD_11595

//ADD_9782 replaced by ADD_11602

//ADD_9781 replaced by ADD_11602

//BasicMUL48_435 replaced by BasicMUL48_970

//BasicMUL48_436 replaced by BasicMUL48_967

//BasicMUL48_437 replaced by BasicMUL48_970

//ADD_9786 replaced by ADD_11602

//ADD_9785 replaced by ADD_11602

//ADD_9784 replaced by ADD_11602

//ADD_9789 replaced by ADD_11601

//ADD_9788 replaced by ADD_11602

//ADD_9787 replaced by ADD_11602

//ADD_9791 replaced by ADD_11602

//ADD_9790 replaced by ADD_11602

//BasicMUL48_438 replaced by BasicMUL48_971

//BasicMUL48_439 replaced by BasicMUL48_970

//BasicMUL48_440 replaced by BasicMUL48_971

//ADD_9794 replaced by ADD_11595

//ADD_9793 replaced by ADD_11602

//ADD_9792 replaced by ADD_11602

//ADD_9797 replaced by ADD_11592

//ADD_9796 replaced by ADD_11602

//ADD_9795 replaced by ADD_11602

//ADD_9800 replaced by ADD_11592

//ADD_9799 replaced by ADD_11602

//ADD_9798 replaced by ADD_11602

//ADD_9803 replaced by ADD_11595

//ADD_9802 replaced by ADD_11602

//ADD_9801 replaced by ADD_11602

//BasicMUL48_441 replaced by BasicMUL48_970

//BasicMUL48_442 replaced by BasicMUL48_967

//BasicMUL48_443 replaced by BasicMUL48_970

//ADD_9806 replaced by ADD_11563

//ADD_9805 replaced by ADD_11602

//ADD_9804 replaced by ADD_11602

//ADD_9809 replaced by ADD_11560

//ADD_9808 replaced by ADD_11602

//ADD_9807 replaced by ADD_11602

//ADD_9812 replaced by ADD_11560

//ADD_9811 replaced by ADD_11602

//ADD_9810 replaced by ADD_11602

//ADD_9815 replaced by ADD_11563

//ADD_9814 replaced by ADD_11602

//ADD_9813 replaced by ADD_11602

//BasicMUL48_444 replaced by BasicMUL48_967

//BasicMUL48_445 replaced by BasicMUL48_958

//BasicMUL48_446 replaced by BasicMUL48_967

//ADD_9818 replaced by ADD_11595

//ADD_9817 replaced by ADD_11602

//ADD_9816 replaced by ADD_11602

//ADD_9821 replaced by ADD_11592

//ADD_9820 replaced by ADD_11602

//ADD_9819 replaced by ADD_11602

//ADD_9824 replaced by ADD_11592

//ADD_9823 replaced by ADD_11602

//ADD_9822 replaced by ADD_11602

//ADD_9827 replaced by ADD_11595

//ADD_9826 replaced by ADD_11602

//ADD_9825 replaced by ADD_11602

//BasicMUL48_447 replaced by BasicMUL48_970

//BasicMUL48_448 replaced by BasicMUL48_967

//BasicMUL48_449 replaced by BasicMUL48_970

//ADD_9830 replaced by ADD_11602

//ADD_9829 replaced by ADD_11602

//ADD_9828 replaced by ADD_11602

//ADD_9833 replaced by ADD_11601

//ADD_9832 replaced by ADD_11602

//ADD_9831 replaced by ADD_11602

//ADD_9835 replaced by ADD_11602

//ADD_9834 replaced by ADD_11602

//BasicMUL48_450 replaced by BasicMUL48_971

//BasicMUL48_451 replaced by BasicMUL48_970

//BasicMUL48_452 replaced by BasicMUL48_971

//ADD_9838 replaced by ADD_11595

//ADD_9837 replaced by ADD_11602

//ADD_9836 replaced by ADD_11602

//ADD_9841 replaced by ADD_11592

//ADD_9840 replaced by ADD_11602

//ADD_9839 replaced by ADD_11602

//ADD_9844 replaced by ADD_11592

//ADD_9843 replaced by ADD_11602

//ADD_9842 replaced by ADD_11602

//ADD_9847 replaced by ADD_11595

//ADD_9846 replaced by ADD_11602

//ADD_9845 replaced by ADD_11602

//BasicMUL48_453 replaced by BasicMUL48_970

//BasicMUL48_454 replaced by BasicMUL48_967

//BasicMUL48_455 replaced by BasicMUL48_970

//ADD_9850 replaced by ADD_11602

//ADD_9849 replaced by ADD_11602

//ADD_9848 replaced by ADD_11602

//ADD_9853 replaced by ADD_11601

//ADD_9852 replaced by ADD_11602

//ADD_9851 replaced by ADD_11602

//ADD_9855 replaced by ADD_11602

//ADD_9854 replaced by ADD_11602

//BasicMUL48_456 replaced by BasicMUL48_971

//BasicMUL48_457 replaced by BasicMUL48_970

//BasicMUL48_458 replaced by BasicMUL48_971

//ADD_9858 replaced by ADD_11602

//ADD_9857 replaced by ADD_11602

//ADD_9856 replaced by ADD_11602

//ADD_9861 replaced by ADD_11601

//ADD_9860 replaced by ADD_11602

//ADD_9859 replaced by ADD_11602

//ADD_9863 replaced by ADD_11602

//ADD_9862 replaced by ADD_11602

//BasicMUL48_459 replaced by BasicMUL48_971

//BasicMUL48_460 replaced by BasicMUL48_970

//BasicMUL48_461 replaced by BasicMUL48_971

//ADD_9866 replaced by ADD_11595

//ADD_9865 replaced by ADD_11602

//ADD_9864 replaced by ADD_11602

//ADD_9869 replaced by ADD_11592

//ADD_9868 replaced by ADD_11602

//ADD_9867 replaced by ADD_11602

//ADD_9872 replaced by ADD_11592

//ADD_9871 replaced by ADD_11602

//ADD_9870 replaced by ADD_11602

//ADD_9875 replaced by ADD_11595

//ADD_9874 replaced by ADD_11602

//ADD_9873 replaced by ADD_11602

//BasicMUL48_462 replaced by BasicMUL48_970

//BasicMUL48_463 replaced by BasicMUL48_967

//BasicMUL48_464 replaced by BasicMUL48_970

//ADD_9878 replaced by ADD_11602

//ADD_9877 replaced by ADD_11602

//ADD_9876 replaced by ADD_11602

//ADD_9881 replaced by ADD_11601

//ADD_9880 replaced by ADD_11602

//ADD_9879 replaced by ADD_11602

//ADD_9883 replaced by ADD_11602

//ADD_9882 replaced by ADD_11602

//BasicMUL48_465 replaced by BasicMUL48_971

//BasicMUL48_466 replaced by BasicMUL48_970

//BasicMUL48_467 replaced by BasicMUL48_971

//ADD_9886 replaced by ADD_11595

//ADD_9885 replaced by ADD_11602

//ADD_9884 replaced by ADD_11602

//ADD_9889 replaced by ADD_11592

//ADD_9888 replaced by ADD_11602

//ADD_9887 replaced by ADD_11602

//ADD_9892 replaced by ADD_11592

//ADD_9891 replaced by ADD_11602

//ADD_9890 replaced by ADD_11602

//ADD_9895 replaced by ADD_11595

//ADD_9894 replaced by ADD_11602

//ADD_9893 replaced by ADD_11602

//BasicMUL48_468 replaced by BasicMUL48_970

//BasicMUL48_469 replaced by BasicMUL48_967

//BasicMUL48_470 replaced by BasicMUL48_970

//ADD_9898 replaced by ADD_11563

//ADD_9897 replaced by ADD_11602

//ADD_9896 replaced by ADD_11602

//ADD_9901 replaced by ADD_11560

//ADD_9900 replaced by ADD_11602

//ADD_9899 replaced by ADD_11602

//ADD_9904 replaced by ADD_11560

//ADD_9903 replaced by ADD_11602

//ADD_9902 replaced by ADD_11602

//ADD_9907 replaced by ADD_11563

//ADD_9906 replaced by ADD_11602

//ADD_9905 replaced by ADD_11602

//BasicMUL48_471 replaced by BasicMUL48_967

//BasicMUL48_472 replaced by BasicMUL48_958

//BasicMUL48_473 replaced by BasicMUL48_967

//ADD_9910 replaced by ADD_11595

//ADD_9909 replaced by ADD_11602

//ADD_9908 replaced by ADD_11602

//ADD_9913 replaced by ADD_11592

//ADD_9912 replaced by ADD_11602

//ADD_9911 replaced by ADD_11602

//ADD_9916 replaced by ADD_11592

//ADD_9915 replaced by ADD_11602

//ADD_9914 replaced by ADD_11602

//ADD_9919 replaced by ADD_11595

//ADD_9918 replaced by ADD_11602

//ADD_9917 replaced by ADD_11602

//BasicMUL48_474 replaced by BasicMUL48_970

//BasicMUL48_475 replaced by BasicMUL48_967

//BasicMUL48_476 replaced by BasicMUL48_970

//ADD_9922 replaced by ADD_11602

//ADD_9921 replaced by ADD_11602

//ADD_9920 replaced by ADD_11602

//ADD_9925 replaced by ADD_11601

//ADD_9924 replaced by ADD_11602

//ADD_9923 replaced by ADD_11602

//ADD_9927 replaced by ADD_11602

//ADD_9926 replaced by ADD_11602

//BasicMUL48_477 replaced by BasicMUL48_971

//BasicMUL48_478 replaced by BasicMUL48_970

//BasicMUL48_479 replaced by BasicMUL48_971

//ADD_9930 replaced by ADD_11595

//ADD_9929 replaced by ADD_11602

//ADD_9928 replaced by ADD_11602

//ADD_9933 replaced by ADD_11592

//ADD_9932 replaced by ADD_11602

//ADD_9931 replaced by ADD_11602

//ADD_9936 replaced by ADD_11592

//ADD_9935 replaced by ADD_11602

//ADD_9934 replaced by ADD_11602

//ADD_9939 replaced by ADD_11595

//ADD_9938 replaced by ADD_11602

//ADD_9937 replaced by ADD_11602

//BasicMUL48_480 replaced by BasicMUL48_970

//BasicMUL48_481 replaced by BasicMUL48_967

//BasicMUL48_482 replaced by BasicMUL48_970

//ADD_9942 replaced by ADD_11602

//ADD_9941 replaced by ADD_11602

//ADD_9940 replaced by ADD_11602

//ADD_9945 replaced by ADD_11601

//ADD_9944 replaced by ADD_11602

//ADD_9943 replaced by ADD_11602

//ADD_9947 replaced by ADD_11602

//ADD_9946 replaced by ADD_11602

//BasicMUL48_483 replaced by BasicMUL48_971

//BasicMUL48_484 replaced by BasicMUL48_970

//BasicMUL48_485 replaced by BasicMUL48_971

//ADD_9950 replaced by ADD_11602

//ADD_9949 replaced by ADD_11602

//ADD_9948 replaced by ADD_11602

//ADD_9953 replaced by ADD_11601

//ADD_9952 replaced by ADD_11602

//ADD_9951 replaced by ADD_11602

//ADD_9955 replaced by ADD_11602

//ADD_9954 replaced by ADD_11602

//BasicMUL48_486 replaced by BasicMUL48_971

//BasicMUL48_487 replaced by BasicMUL48_970

//BasicMUL48_488 replaced by BasicMUL48_971

//ADD_9958 replaced by ADD_11595

//ADD_9957 replaced by ADD_11602

//ADD_9956 replaced by ADD_11602

//ADD_9961 replaced by ADD_11592

//ADD_9960 replaced by ADD_11602

//ADD_9959 replaced by ADD_11602

//ADD_9964 replaced by ADD_11592

//ADD_9963 replaced by ADD_11602

//ADD_9962 replaced by ADD_11602

//ADD_9967 replaced by ADD_11595

//ADD_9966 replaced by ADD_11602

//ADD_9965 replaced by ADD_11602

//BasicMUL48_489 replaced by BasicMUL48_970

//BasicMUL48_490 replaced by BasicMUL48_967

//BasicMUL48_491 replaced by BasicMUL48_970

//ADD_9970 replaced by ADD_11602

//ADD_9969 replaced by ADD_11602

//ADD_9968 replaced by ADD_11602

//ADD_9973 replaced by ADD_11601

//ADD_9972 replaced by ADD_11602

//ADD_9971 replaced by ADD_11602

//ADD_9975 replaced by ADD_11602

//ADD_9974 replaced by ADD_11602

//BasicMUL48_492 replaced by BasicMUL48_971

//BasicMUL48_493 replaced by BasicMUL48_970

//BasicMUL48_494 replaced by BasicMUL48_971

//ADD_9978 replaced by ADD_11595

//ADD_9977 replaced by ADD_11602

//ADD_9976 replaced by ADD_11602

//ADD_9981 replaced by ADD_11592

//ADD_9980 replaced by ADD_11602

//ADD_9979 replaced by ADD_11602

//ADD_9984 replaced by ADD_11592

//ADD_9983 replaced by ADD_11602

//ADD_9982 replaced by ADD_11602

//ADD_9987 replaced by ADD_11595

//ADD_9986 replaced by ADD_11602

//ADD_9985 replaced by ADD_11602

//BasicMUL48_495 replaced by BasicMUL48_970

//BasicMUL48_496 replaced by BasicMUL48_967

//BasicMUL48_497 replaced by BasicMUL48_970

//ADD_9990 replaced by ADD_11563

//ADD_9989 replaced by ADD_11602

//ADD_9988 replaced by ADD_11602

//ADD_9993 replaced by ADD_11560

//ADD_9992 replaced by ADD_11602

//ADD_9991 replaced by ADD_11602

//ADD_9996 replaced by ADD_11560

//ADD_9995 replaced by ADD_11602

//ADD_9994 replaced by ADD_11602

//ADD_9999 replaced by ADD_11563

//ADD_9998 replaced by ADD_11602

//ADD_9997 replaced by ADD_11602

//BasicMUL48_498 replaced by BasicMUL48_967

//BasicMUL48_499 replaced by BasicMUL48_958

//BasicMUL48_500 replaced by BasicMUL48_967

//ADD_10002 replaced by ADD_11595

//ADD_10001 replaced by ADD_11602

//ADD_10000 replaced by ADD_11602

//ADD_10005 replaced by ADD_11592

//ADD_10004 replaced by ADD_11602

//ADD_10003 replaced by ADD_11602

//ADD_10008 replaced by ADD_11592

//ADD_10007 replaced by ADD_11602

//ADD_10006 replaced by ADD_11602

//ADD_10011 replaced by ADD_11595

//ADD_10010 replaced by ADD_11602

//ADD_10009 replaced by ADD_11602

//BasicMUL48_501 replaced by BasicMUL48_970

//BasicMUL48_502 replaced by BasicMUL48_967

//BasicMUL48_503 replaced by BasicMUL48_970

//ADD_10014 replaced by ADD_11602

//ADD_10013 replaced by ADD_11602

//ADD_10012 replaced by ADD_11602

//ADD_10017 replaced by ADD_11601

//ADD_10016 replaced by ADD_11602

//ADD_10015 replaced by ADD_11602

//ADD_10019 replaced by ADD_11602

//ADD_10018 replaced by ADD_11602

//BasicMUL48_504 replaced by BasicMUL48_971

//BasicMUL48_505 replaced by BasicMUL48_970

//BasicMUL48_506 replaced by BasicMUL48_971

//ADD_10022 replaced by ADD_11595

//ADD_10021 replaced by ADD_11602

//ADD_10020 replaced by ADD_11602

//ADD_10025 replaced by ADD_11592

//ADD_10024 replaced by ADD_11602

//ADD_10023 replaced by ADD_11602

//ADD_10028 replaced by ADD_11592

//ADD_10027 replaced by ADD_11602

//ADD_10026 replaced by ADD_11602

//ADD_10031 replaced by ADD_11595

//ADD_10030 replaced by ADD_11602

//ADD_10029 replaced by ADD_11602

//BasicMUL48_507 replaced by BasicMUL48_970

//BasicMUL48_508 replaced by BasicMUL48_967

//BasicMUL48_509 replaced by BasicMUL48_970

//ADD_10034 replaced by ADD_11602

//ADD_10033 replaced by ADD_11602

//ADD_10032 replaced by ADD_11602

//ADD_10037 replaced by ADD_11601

//ADD_10036 replaced by ADD_11602

//ADD_10035 replaced by ADD_11602

//ADD_10039 replaced by ADD_11602

//ADD_10038 replaced by ADD_11602

//BasicMUL48_510 replaced by BasicMUL48_971

//BasicMUL48_511 replaced by BasicMUL48_970

//BasicMUL48_512 replaced by BasicMUL48_971

//ADD_10042 replaced by ADD_11602

//ADD_10041 replaced by ADD_11602

//ADD_10040 replaced by ADD_11602

//ADD_10045 replaced by ADD_11601

//ADD_10044 replaced by ADD_11602

//ADD_10043 replaced by ADD_11602

//ADD_10047 replaced by ADD_11602

//ADD_10046 replaced by ADD_11602

//BasicMUL48_513 replaced by BasicMUL48_971

//BasicMUL48_514 replaced by BasicMUL48_970

//BasicMUL48_515 replaced by BasicMUL48_971

//ADD_10050 replaced by ADD_11595

//ADD_10049 replaced by ADD_11602

//ADD_10048 replaced by ADD_11602

//ADD_10053 replaced by ADD_11592

//ADD_10052 replaced by ADD_11602

//ADD_10051 replaced by ADD_11602

//ADD_10056 replaced by ADD_11592

//ADD_10055 replaced by ADD_11602

//ADD_10054 replaced by ADD_11602

//ADD_10059 replaced by ADD_11595

//ADD_10058 replaced by ADD_11602

//ADD_10057 replaced by ADD_11602

//BasicMUL48_516 replaced by BasicMUL48_970

//BasicMUL48_517 replaced by BasicMUL48_967

//BasicMUL48_518 replaced by BasicMUL48_970

//ADD_10062 replaced by ADD_11602

//ADD_10061 replaced by ADD_11602

//ADD_10060 replaced by ADD_11602

//ADD_10065 replaced by ADD_11601

//ADD_10064 replaced by ADD_11602

//ADD_10063 replaced by ADD_11602

//ADD_10067 replaced by ADD_11602

//ADD_10066 replaced by ADD_11602

//BasicMUL48_519 replaced by BasicMUL48_971

//BasicMUL48_520 replaced by BasicMUL48_970

//BasicMUL48_521 replaced by BasicMUL48_971

//ADD_10070 replaced by ADD_11595

//ADD_10069 replaced by ADD_11602

//ADD_10068 replaced by ADD_11602

//ADD_10073 replaced by ADD_11592

//ADD_10072 replaced by ADD_11602

//ADD_10071 replaced by ADD_11602

//ADD_10076 replaced by ADD_11592

//ADD_10075 replaced by ADD_11602

//ADD_10074 replaced by ADD_11602

//ADD_10079 replaced by ADD_11595

//ADD_10078 replaced by ADD_11602

//ADD_10077 replaced by ADD_11602

//BasicMUL48_522 replaced by BasicMUL48_970

//BasicMUL48_523 replaced by BasicMUL48_967

//BasicMUL48_524 replaced by BasicMUL48_970

//ADD_10082 replaced by ADD_11563

//ADD_10081 replaced by ADD_11602

//ADD_10080 replaced by ADD_11602

//ADD_10085 replaced by ADD_11560

//ADD_10084 replaced by ADD_11602

//ADD_10083 replaced by ADD_11602

//ADD_10088 replaced by ADD_11560

//ADD_10087 replaced by ADD_11602

//ADD_10086 replaced by ADD_11602

//ADD_10091 replaced by ADD_11563

//ADD_10090 replaced by ADD_11602

//ADD_10089 replaced by ADD_11602

//BasicMUL48_525 replaced by BasicMUL48_967

//BasicMUL48_526 replaced by BasicMUL48_958

//BasicMUL48_527 replaced by BasicMUL48_967

//ADD_10094 replaced by ADD_11595

//ADD_10093 replaced by ADD_11602

//ADD_10092 replaced by ADD_11602

//ADD_10097 replaced by ADD_11592

//ADD_10096 replaced by ADD_11602

//ADD_10095 replaced by ADD_11602

//ADD_10100 replaced by ADD_11592

//ADD_10099 replaced by ADD_11602

//ADD_10098 replaced by ADD_11602

//ADD_10103 replaced by ADD_11595

//ADD_10102 replaced by ADD_11602

//ADD_10101 replaced by ADD_11602

//BasicMUL48_528 replaced by BasicMUL48_970

//BasicMUL48_529 replaced by BasicMUL48_967

//BasicMUL48_530 replaced by BasicMUL48_970

//ADD_10106 replaced by ADD_11602

//ADD_10105 replaced by ADD_11602

//ADD_10104 replaced by ADD_11602

//ADD_10109 replaced by ADD_11601

//ADD_10108 replaced by ADD_11602

//ADD_10107 replaced by ADD_11602

//ADD_10111 replaced by ADD_11602

//ADD_10110 replaced by ADD_11602

//BasicMUL48_531 replaced by BasicMUL48_971

//BasicMUL48_532 replaced by BasicMUL48_970

//BasicMUL48_533 replaced by BasicMUL48_971

//ADD_10114 replaced by ADD_11595

//ADD_10113 replaced by ADD_11602

//ADD_10112 replaced by ADD_11602

//ADD_10117 replaced by ADD_11592

//ADD_10116 replaced by ADD_11602

//ADD_10115 replaced by ADD_11602

//ADD_10120 replaced by ADD_11592

//ADD_10119 replaced by ADD_11602

//ADD_10118 replaced by ADD_11602

//ADD_10123 replaced by ADD_11595

//ADD_10122 replaced by ADD_11602

//ADD_10121 replaced by ADD_11602

//BasicMUL48_534 replaced by BasicMUL48_970

//BasicMUL48_535 replaced by BasicMUL48_967

//BasicMUL48_536 replaced by BasicMUL48_970

//ADD_10126 replaced by ADD_11602

//ADD_10125 replaced by ADD_11602

//ADD_10124 replaced by ADD_11602

//ADD_10129 replaced by ADD_11601

//ADD_10128 replaced by ADD_11602

//ADD_10127 replaced by ADD_11602

//ADD_10131 replaced by ADD_11602

//ADD_10130 replaced by ADD_11602

//BasicMUL48_537 replaced by BasicMUL48_971

//BasicMUL48_538 replaced by BasicMUL48_970

//BasicMUL48_539 replaced by BasicMUL48_971

//ADD_10134 replaced by ADD_11602

//ADD_10133 replaced by ADD_11602

//ADD_10132 replaced by ADD_11602

//ADD_10137 replaced by ADD_11601

//ADD_10136 replaced by ADD_11602

//ADD_10135 replaced by ADD_11602

//ADD_10139 replaced by ADD_11602

//ADD_10138 replaced by ADD_11602

//BasicMUL48_540 replaced by BasicMUL48_971

//BasicMUL48_541 replaced by BasicMUL48_970

//BasicMUL48_542 replaced by BasicMUL48_971

//ADD_10142 replaced by ADD_11595

//ADD_10141 replaced by ADD_11602

//ADD_10140 replaced by ADD_11602

//ADD_10145 replaced by ADD_11592

//ADD_10144 replaced by ADD_11602

//ADD_10143 replaced by ADD_11602

//ADD_10148 replaced by ADD_11592

//ADD_10147 replaced by ADD_11602

//ADD_10146 replaced by ADD_11602

//ADD_10151 replaced by ADD_11595

//ADD_10150 replaced by ADD_11602

//ADD_10149 replaced by ADD_11602

//BasicMUL48_543 replaced by BasicMUL48_970

//BasicMUL48_544 replaced by BasicMUL48_967

//BasicMUL48_545 replaced by BasicMUL48_970

//ADD_10154 replaced by ADD_11602

//ADD_10153 replaced by ADD_11602

//ADD_10152 replaced by ADD_11602

//ADD_10157 replaced by ADD_11601

//ADD_10156 replaced by ADD_11602

//ADD_10155 replaced by ADD_11602

//ADD_10159 replaced by ADD_11602

//ADD_10158 replaced by ADD_11602

//BasicMUL48_546 replaced by BasicMUL48_971

//BasicMUL48_547 replaced by BasicMUL48_970

//BasicMUL48_548 replaced by BasicMUL48_971

//ADD_10162 replaced by ADD_11595

//ADD_10161 replaced by ADD_11602

//ADD_10160 replaced by ADD_11602

//ADD_10165 replaced by ADD_11592

//ADD_10164 replaced by ADD_11602

//ADD_10163 replaced by ADD_11602

//ADD_10168 replaced by ADD_11592

//ADD_10167 replaced by ADD_11602

//ADD_10166 replaced by ADD_11602

//ADD_10171 replaced by ADD_11595

//ADD_10170 replaced by ADD_11602

//ADD_10169 replaced by ADD_11602

//BasicMUL48_549 replaced by BasicMUL48_970

//BasicMUL48_550 replaced by BasicMUL48_967

//BasicMUL48_551 replaced by BasicMUL48_970

//ADD_10174 replaced by ADD_11563

//ADD_10173 replaced by ADD_11602

//ADD_10172 replaced by ADD_11602

//ADD_10177 replaced by ADD_11560

//ADD_10176 replaced by ADD_11602

//ADD_10175 replaced by ADD_11602

//ADD_10180 replaced by ADD_11560

//ADD_10179 replaced by ADD_11602

//ADD_10178 replaced by ADD_11602

//ADD_10183 replaced by ADD_11563

//ADD_10182 replaced by ADD_11602

//ADD_10181 replaced by ADD_11602

//BasicMUL48_552 replaced by BasicMUL48_967

//BasicMUL48_553 replaced by BasicMUL48_958

//BasicMUL48_554 replaced by BasicMUL48_967

//ADD_10186 replaced by ADD_11595

//ADD_10185 replaced by ADD_11602

//ADD_10184 replaced by ADD_11602

//ADD_10189 replaced by ADD_11592

//ADD_10188 replaced by ADD_11602

//ADD_10187 replaced by ADD_11602

//ADD_10192 replaced by ADD_11592

//ADD_10191 replaced by ADD_11602

//ADD_10190 replaced by ADD_11602

//ADD_10195 replaced by ADD_11595

//ADD_10194 replaced by ADD_11602

//ADD_10193 replaced by ADD_11602

//BasicMUL48_555 replaced by BasicMUL48_970

//BasicMUL48_556 replaced by BasicMUL48_967

//BasicMUL48_557 replaced by BasicMUL48_970

//ADD_10198 replaced by ADD_11602

//ADD_10197 replaced by ADD_11602

//ADD_10196 replaced by ADD_11602

//ADD_10201 replaced by ADD_11601

//ADD_10200 replaced by ADD_11602

//ADD_10199 replaced by ADD_11602

//ADD_10203 replaced by ADD_11602

//ADD_10202 replaced by ADD_11602

//BasicMUL48_558 replaced by BasicMUL48_971

//BasicMUL48_559 replaced by BasicMUL48_970

//BasicMUL48_560 replaced by BasicMUL48_971

//ADD_10206 replaced by ADD_11595

//ADD_10205 replaced by ADD_11602

//ADD_10204 replaced by ADD_11602

//ADD_10209 replaced by ADD_11592

//ADD_10208 replaced by ADD_11602

//ADD_10207 replaced by ADD_11602

//ADD_10212 replaced by ADD_11592

//ADD_10211 replaced by ADD_11602

//ADD_10210 replaced by ADD_11602

//ADD_10215 replaced by ADD_11595

//ADD_10214 replaced by ADD_11602

//ADD_10213 replaced by ADD_11602

//BasicMUL48_561 replaced by BasicMUL48_970

//BasicMUL48_562 replaced by BasicMUL48_967

//BasicMUL48_563 replaced by BasicMUL48_970

//ADD_10218 replaced by ADD_11602

//ADD_10217 replaced by ADD_11602

//ADD_10216 replaced by ADD_11602

//ADD_10221 replaced by ADD_11601

//ADD_10220 replaced by ADD_11602

//ADD_10219 replaced by ADD_11602

//ADD_10223 replaced by ADD_11602

//ADD_10222 replaced by ADD_11602

//BasicMUL48_564 replaced by BasicMUL48_971

//BasicMUL48_565 replaced by BasicMUL48_970

//BasicMUL48_566 replaced by BasicMUL48_971

//ADD_10226 replaced by ADD_11602

//ADD_10225 replaced by ADD_11602

//ADD_10224 replaced by ADD_11602

//ADD_10229 replaced by ADD_11601

//ADD_10228 replaced by ADD_11602

//ADD_10227 replaced by ADD_11602

//ADD_10231 replaced by ADD_11602

//ADD_10230 replaced by ADD_11602

//BasicMUL48_567 replaced by BasicMUL48_971

//BasicMUL48_568 replaced by BasicMUL48_970

//BasicMUL48_569 replaced by BasicMUL48_971

//ADD_10234 replaced by ADD_11595

//ADD_10233 replaced by ADD_11602

//ADD_10232 replaced by ADD_11602

//ADD_10237 replaced by ADD_11592

//ADD_10236 replaced by ADD_11602

//ADD_10235 replaced by ADD_11602

//ADD_10240 replaced by ADD_11592

//ADD_10239 replaced by ADD_11602

//ADD_10238 replaced by ADD_11602

//ADD_10243 replaced by ADD_11595

//ADD_10242 replaced by ADD_11602

//ADD_10241 replaced by ADD_11602

//BasicMUL48_570 replaced by BasicMUL48_970

//BasicMUL48_571 replaced by BasicMUL48_967

//BasicMUL48_572 replaced by BasicMUL48_970

//ADD_10246 replaced by ADD_11602

//ADD_10245 replaced by ADD_11602

//ADD_10244 replaced by ADD_11602

//ADD_10249 replaced by ADD_11601

//ADD_10248 replaced by ADD_11602

//ADD_10247 replaced by ADD_11602

//ADD_10251 replaced by ADD_11602

//ADD_10250 replaced by ADD_11602

//BasicMUL48_573 replaced by BasicMUL48_971

//BasicMUL48_574 replaced by BasicMUL48_970

//BasicMUL48_575 replaced by BasicMUL48_971

//ADD_10254 replaced by ADD_11595

//ADD_10253 replaced by ADD_11602

//ADD_10252 replaced by ADD_11602

//ADD_10257 replaced by ADD_11592

//ADD_10256 replaced by ADD_11602

//ADD_10255 replaced by ADD_11602

//ADD_10260 replaced by ADD_11592

//ADD_10259 replaced by ADD_11602

//ADD_10258 replaced by ADD_11602

//ADD_10263 replaced by ADD_11595

//ADD_10262 replaced by ADD_11602

//ADD_10261 replaced by ADD_11602

//BasicMUL48_576 replaced by BasicMUL48_970

//BasicMUL48_577 replaced by BasicMUL48_967

//BasicMUL48_578 replaced by BasicMUL48_970

//ADD_10266 replaced by ADD_11563

//ADD_10265 replaced by ADD_11602

//ADD_10264 replaced by ADD_11602

//ADD_10269 replaced by ADD_11560

//ADD_10268 replaced by ADD_11602

//ADD_10267 replaced by ADD_11602

//ADD_10272 replaced by ADD_11560

//ADD_10271 replaced by ADD_11602

//ADD_10270 replaced by ADD_11602

//ADD_10275 replaced by ADD_11563

//ADD_10274 replaced by ADD_11602

//ADD_10273 replaced by ADD_11602

//BasicMUL48_579 replaced by BasicMUL48_967

//BasicMUL48_580 replaced by BasicMUL48_958

//BasicMUL48_581 replaced by BasicMUL48_967

//ADD_10278 replaced by ADD_11595

//ADD_10277 replaced by ADD_11602

//ADD_10276 replaced by ADD_11602

//ADD_10281 replaced by ADD_11592

//ADD_10280 replaced by ADD_11602

//ADD_10279 replaced by ADD_11602

//ADD_10284 replaced by ADD_11592

//ADD_10283 replaced by ADD_11602

//ADD_10282 replaced by ADD_11602

//ADD_10287 replaced by ADD_11595

//ADD_10286 replaced by ADD_11602

//ADD_10285 replaced by ADD_11602

//BasicMUL48_582 replaced by BasicMUL48_970

//BasicMUL48_583 replaced by BasicMUL48_967

//BasicMUL48_584 replaced by BasicMUL48_970

//ADD_10290 replaced by ADD_11602

//ADD_10289 replaced by ADD_11602

//ADD_10288 replaced by ADD_11602

//ADD_10293 replaced by ADD_11601

//ADD_10292 replaced by ADD_11602

//ADD_10291 replaced by ADD_11602

//ADD_10295 replaced by ADD_11602

//ADD_10294 replaced by ADD_11602

//BasicMUL48_585 replaced by BasicMUL48_971

//BasicMUL48_586 replaced by BasicMUL48_970

//BasicMUL48_587 replaced by BasicMUL48_971

//ADD_10298 replaced by ADD_11595

//ADD_10297 replaced by ADD_11602

//ADD_10296 replaced by ADD_11602

//ADD_10301 replaced by ADD_11592

//ADD_10300 replaced by ADD_11602

//ADD_10299 replaced by ADD_11602

//ADD_10304 replaced by ADD_11592

//ADD_10303 replaced by ADD_11602

//ADD_10302 replaced by ADD_11602

//ADD_10307 replaced by ADD_11595

//ADD_10306 replaced by ADD_11602

//ADD_10305 replaced by ADD_11602

//BasicMUL48_588 replaced by BasicMUL48_970

//BasicMUL48_589 replaced by BasicMUL48_967

//BasicMUL48_590 replaced by BasicMUL48_970

//ADD_10310 replaced by ADD_11602

//ADD_10309 replaced by ADD_11602

//ADD_10308 replaced by ADD_11602

//ADD_10313 replaced by ADD_11601

//ADD_10312 replaced by ADD_11602

//ADD_10311 replaced by ADD_11602

//ADD_10315 replaced by ADD_11602

//ADD_10314 replaced by ADD_11602

//BasicMUL48_591 replaced by BasicMUL48_971

//BasicMUL48_592 replaced by BasicMUL48_970

//BasicMUL48_593 replaced by BasicMUL48_971

//ADD_10318 replaced by ADD_11602

//ADD_10317 replaced by ADD_11602

//ADD_10316 replaced by ADD_11602

//ADD_10321 replaced by ADD_11601

//ADD_10320 replaced by ADD_11602

//ADD_10319 replaced by ADD_11602

//ADD_10323 replaced by ADD_11602

//ADD_10322 replaced by ADD_11602

//BasicMUL48_594 replaced by BasicMUL48_971

//BasicMUL48_595 replaced by BasicMUL48_970

//BasicMUL48_596 replaced by BasicMUL48_971

//ADD_10326 replaced by ADD_11595

//ADD_10325 replaced by ADD_11602

//ADD_10324 replaced by ADD_11602

//ADD_10329 replaced by ADD_11592

//ADD_10328 replaced by ADD_11602

//ADD_10327 replaced by ADD_11602

//ADD_10332 replaced by ADD_11592

//ADD_10331 replaced by ADD_11602

//ADD_10330 replaced by ADD_11602

//ADD_10335 replaced by ADD_11595

//ADD_10334 replaced by ADD_11602

//ADD_10333 replaced by ADD_11602

//BasicMUL48_597 replaced by BasicMUL48_970

//BasicMUL48_598 replaced by BasicMUL48_967

//BasicMUL48_599 replaced by BasicMUL48_970

//ADD_10338 replaced by ADD_11602

//ADD_10337 replaced by ADD_11602

//ADD_10336 replaced by ADD_11602

//ADD_10341 replaced by ADD_11601

//ADD_10340 replaced by ADD_11602

//ADD_10339 replaced by ADD_11602

//ADD_10343 replaced by ADD_11602

//ADD_10342 replaced by ADD_11602

//BasicMUL48_600 replaced by BasicMUL48_971

//BasicMUL48_601 replaced by BasicMUL48_970

//BasicMUL48_602 replaced by BasicMUL48_971

//ADD_10346 replaced by ADD_11595

//ADD_10345 replaced by ADD_11602

//ADD_10344 replaced by ADD_11602

//ADD_10349 replaced by ADD_11592

//ADD_10348 replaced by ADD_11602

//ADD_10347 replaced by ADD_11602

//ADD_10352 replaced by ADD_11592

//ADD_10351 replaced by ADD_11602

//ADD_10350 replaced by ADD_11602

//ADD_10355 replaced by ADD_11595

//ADD_10354 replaced by ADD_11602

//ADD_10353 replaced by ADD_11602

//BasicMUL48_603 replaced by BasicMUL48_970

//BasicMUL48_604 replaced by BasicMUL48_967

//BasicMUL48_605 replaced by BasicMUL48_970

//ADD_10358 replaced by ADD_11563

//ADD_10357 replaced by ADD_11602

//ADD_10356 replaced by ADD_11602

//ADD_10361 replaced by ADD_11560

//ADD_10360 replaced by ADD_11602

//ADD_10359 replaced by ADD_11602

//ADD_10364 replaced by ADD_11560

//ADD_10363 replaced by ADD_11602

//ADD_10362 replaced by ADD_11602

//ADD_10367 replaced by ADD_11563

//ADD_10366 replaced by ADD_11602

//ADD_10365 replaced by ADD_11602

//BasicMUL48_606 replaced by BasicMUL48_967

//BasicMUL48_607 replaced by BasicMUL48_958

//BasicMUL48_608 replaced by BasicMUL48_967

//ADD_10370 replaced by ADD_11595

//ADD_10369 replaced by ADD_11602

//ADD_10368 replaced by ADD_11602

//ADD_10373 replaced by ADD_11592

//ADD_10372 replaced by ADD_11602

//ADD_10371 replaced by ADD_11602

//ADD_10376 replaced by ADD_11592

//ADD_10375 replaced by ADD_11602

//ADD_10374 replaced by ADD_11602

//ADD_10379 replaced by ADD_11595

//ADD_10378 replaced by ADD_11602

//ADD_10377 replaced by ADD_11602

//BasicMUL48_609 replaced by BasicMUL48_970

//BasicMUL48_610 replaced by BasicMUL48_967

//BasicMUL48_611 replaced by BasicMUL48_970

//ADD_10382 replaced by ADD_11602

//ADD_10381 replaced by ADD_11602

//ADD_10380 replaced by ADD_11602

//ADD_10385 replaced by ADD_11601

//ADD_10384 replaced by ADD_11602

//ADD_10383 replaced by ADD_11602

//ADD_10387 replaced by ADD_11602

//ADD_10386 replaced by ADD_11602

//BasicMUL48_612 replaced by BasicMUL48_971

//BasicMUL48_613 replaced by BasicMUL48_970

//BasicMUL48_614 replaced by BasicMUL48_971

//ADD_10390 replaced by ADD_11595

//ADD_10389 replaced by ADD_11602

//ADD_10388 replaced by ADD_11602

//ADD_10393 replaced by ADD_11592

//ADD_10392 replaced by ADD_11602

//ADD_10391 replaced by ADD_11602

//ADD_10396 replaced by ADD_11592

//ADD_10395 replaced by ADD_11602

//ADD_10394 replaced by ADD_11602

//ADD_10399 replaced by ADD_11595

//ADD_10398 replaced by ADD_11602

//ADD_10397 replaced by ADD_11602

//BasicMUL48_615 replaced by BasicMUL48_970

//BasicMUL48_616 replaced by BasicMUL48_967

//BasicMUL48_617 replaced by BasicMUL48_970

//ADD_10402 replaced by ADD_11602

//ADD_10401 replaced by ADD_11602

//ADD_10400 replaced by ADD_11602

//ADD_10405 replaced by ADD_11601

//ADD_10404 replaced by ADD_11602

//ADD_10403 replaced by ADD_11602

//ADD_10407 replaced by ADD_11602

//ADD_10406 replaced by ADD_11602

//BasicMUL48_618 replaced by BasicMUL48_971

//BasicMUL48_619 replaced by BasicMUL48_970

//BasicMUL48_620 replaced by BasicMUL48_971

//ADD_10410 replaced by ADD_11602

//ADD_10409 replaced by ADD_11602

//ADD_10408 replaced by ADD_11602

//ADD_10413 replaced by ADD_11601

//ADD_10412 replaced by ADD_11602

//ADD_10411 replaced by ADD_11602

//ADD_10415 replaced by ADD_11602

//ADD_10414 replaced by ADD_11602

//BasicMUL48_621 replaced by BasicMUL48_971

//BasicMUL48_622 replaced by BasicMUL48_970

//BasicMUL48_623 replaced by BasicMUL48_971

//ADD_10418 replaced by ADD_11595

//ADD_10417 replaced by ADD_11602

//ADD_10416 replaced by ADD_11602

//ADD_10421 replaced by ADD_11592

//ADD_10420 replaced by ADD_11602

//ADD_10419 replaced by ADD_11602

//ADD_10424 replaced by ADD_11592

//ADD_10423 replaced by ADD_11602

//ADD_10422 replaced by ADD_11602

//ADD_10427 replaced by ADD_11595

//ADD_10426 replaced by ADD_11602

//ADD_10425 replaced by ADD_11602

//BasicMUL48_624 replaced by BasicMUL48_970

//BasicMUL48_625 replaced by BasicMUL48_967

//BasicMUL48_626 replaced by BasicMUL48_970

//ADD_10430 replaced by ADD_11602

//ADD_10429 replaced by ADD_11602

//ADD_10428 replaced by ADD_11602

//ADD_10433 replaced by ADD_11601

//ADD_10432 replaced by ADD_11602

//ADD_10431 replaced by ADD_11602

//ADD_10435 replaced by ADD_11602

//ADD_10434 replaced by ADD_11602

//BasicMUL48_627 replaced by BasicMUL48_971

//BasicMUL48_628 replaced by BasicMUL48_970

//BasicMUL48_629 replaced by BasicMUL48_971

//ADD_10438 replaced by ADD_11595

//ADD_10437 replaced by ADD_11602

//ADD_10436 replaced by ADD_11602

//ADD_10441 replaced by ADD_11592

//ADD_10440 replaced by ADD_11602

//ADD_10439 replaced by ADD_11602

//ADD_10444 replaced by ADD_11592

//ADD_10443 replaced by ADD_11602

//ADD_10442 replaced by ADD_11602

//ADD_10447 replaced by ADD_11595

//ADD_10446 replaced by ADD_11602

//ADD_10445 replaced by ADD_11602

//BasicMUL48_630 replaced by BasicMUL48_970

//BasicMUL48_631 replaced by BasicMUL48_967

//BasicMUL48_632 replaced by BasicMUL48_970

//ADD_10450 replaced by ADD_11563

//ADD_10449 replaced by ADD_11602

//ADD_10448 replaced by ADD_11602

//ADD_10453 replaced by ADD_11560

//ADD_10452 replaced by ADD_11602

//ADD_10451 replaced by ADD_11602

//ADD_10456 replaced by ADD_11560

//ADD_10455 replaced by ADD_11602

//ADD_10454 replaced by ADD_11602

//ADD_10459 replaced by ADD_11563

//ADD_10458 replaced by ADD_11602

//ADD_10457 replaced by ADD_11602

//BasicMUL48_633 replaced by BasicMUL48_967

//BasicMUL48_634 replaced by BasicMUL48_958

//BasicMUL48_635 replaced by BasicMUL48_967

//ADD_10462 replaced by ADD_11595

//ADD_10461 replaced by ADD_11602

//ADD_10460 replaced by ADD_11602

//ADD_10465 replaced by ADD_11592

//ADD_10464 replaced by ADD_11602

//ADD_10463 replaced by ADD_11602

//ADD_10468 replaced by ADD_11592

//ADD_10467 replaced by ADD_11602

//ADD_10466 replaced by ADD_11602

//ADD_10471 replaced by ADD_11595

//ADD_10470 replaced by ADD_11602

//ADD_10469 replaced by ADD_11602

//BasicMUL48_636 replaced by BasicMUL48_970

//BasicMUL48_637 replaced by BasicMUL48_967

//BasicMUL48_638 replaced by BasicMUL48_970

//ADD_10474 replaced by ADD_11602

//ADD_10473 replaced by ADD_11602

//ADD_10472 replaced by ADD_11602

//ADD_10477 replaced by ADD_11601

//ADD_10476 replaced by ADD_11602

//ADD_10475 replaced by ADD_11602

//ADD_10479 replaced by ADD_11602

//ADD_10478 replaced by ADD_11602

//BasicMUL48_639 replaced by BasicMUL48_971

//BasicMUL48_640 replaced by BasicMUL48_970

//BasicMUL48_641 replaced by BasicMUL48_971

//ADD_10482 replaced by ADD_11595

//ADD_10481 replaced by ADD_11602

//ADD_10480 replaced by ADD_11602

//ADD_10485 replaced by ADD_11592

//ADD_10484 replaced by ADD_11602

//ADD_10483 replaced by ADD_11602

//ADD_10488 replaced by ADD_11592

//ADD_10487 replaced by ADD_11602

//ADD_10486 replaced by ADD_11602

//ADD_10491 replaced by ADD_11595

//ADD_10490 replaced by ADD_11602

//ADD_10489 replaced by ADD_11602

//BasicMUL48_642 replaced by BasicMUL48_970

//BasicMUL48_643 replaced by BasicMUL48_967

//BasicMUL48_644 replaced by BasicMUL48_970

//ADD_10494 replaced by ADD_11602

//ADD_10493 replaced by ADD_11602

//ADD_10492 replaced by ADD_11602

//ADD_10497 replaced by ADD_11601

//ADD_10496 replaced by ADD_11602

//ADD_10495 replaced by ADD_11602

//ADD_10499 replaced by ADD_11602

//ADD_10498 replaced by ADD_11602

//BasicMUL48_645 replaced by BasicMUL48_971

//BasicMUL48_646 replaced by BasicMUL48_970

//BasicMUL48_647 replaced by BasicMUL48_971

//ADD_10502 replaced by ADD_11602

//ADD_10501 replaced by ADD_11602

//ADD_10500 replaced by ADD_11602

//ADD_10505 replaced by ADD_11601

//ADD_10504 replaced by ADD_11602

//ADD_10503 replaced by ADD_11602

//ADD_10507 replaced by ADD_11602

//ADD_10506 replaced by ADD_11602

//BasicMUL48_648 replaced by BasicMUL48_971

//BasicMUL48_649 replaced by BasicMUL48_970

//BasicMUL48_650 replaced by BasicMUL48_971

//ADD_10510 replaced by ADD_11595

//ADD_10509 replaced by ADD_11602

//ADD_10508 replaced by ADD_11602

//ADD_10513 replaced by ADD_11592

//ADD_10512 replaced by ADD_11602

//ADD_10511 replaced by ADD_11602

//ADD_10516 replaced by ADD_11592

//ADD_10515 replaced by ADD_11602

//ADD_10514 replaced by ADD_11602

//ADD_10519 replaced by ADD_11595

//ADD_10518 replaced by ADD_11602

//ADD_10517 replaced by ADD_11602

//BasicMUL48_651 replaced by BasicMUL48_970

//BasicMUL48_652 replaced by BasicMUL48_967

//BasicMUL48_653 replaced by BasicMUL48_970

//ADD_10522 replaced by ADD_11602

//ADD_10521 replaced by ADD_11602

//ADD_10520 replaced by ADD_11602

//ADD_10525 replaced by ADD_11601

//ADD_10524 replaced by ADD_11602

//ADD_10523 replaced by ADD_11602

//ADD_10527 replaced by ADD_11602

//ADD_10526 replaced by ADD_11602

//BasicMUL48_654 replaced by BasicMUL48_971

//BasicMUL48_655 replaced by BasicMUL48_970

//BasicMUL48_656 replaced by BasicMUL48_971

//ADD_10530 replaced by ADD_11595

//ADD_10529 replaced by ADD_11602

//ADD_10528 replaced by ADD_11602

//ADD_10533 replaced by ADD_11592

//ADD_10532 replaced by ADD_11602

//ADD_10531 replaced by ADD_11602

//ADD_10536 replaced by ADD_11592

//ADD_10535 replaced by ADD_11602

//ADD_10534 replaced by ADD_11602

//ADD_10539 replaced by ADD_11595

//ADD_10538 replaced by ADD_11602

//ADD_10537 replaced by ADD_11602

//BasicMUL48_657 replaced by BasicMUL48_970

//BasicMUL48_658 replaced by BasicMUL48_967

//BasicMUL48_659 replaced by BasicMUL48_970

//ADD_10542 replaced by ADD_11563

//ADD_10541 replaced by ADD_11602

//ADD_10540 replaced by ADD_11602

//ADD_10545 replaced by ADD_11560

//ADD_10544 replaced by ADD_11602

//ADD_10543 replaced by ADD_11602

//ADD_10548 replaced by ADD_11560

//ADD_10547 replaced by ADD_11602

//ADD_10546 replaced by ADD_11602

//ADD_10551 replaced by ADD_11563

//ADD_10550 replaced by ADD_11602

//ADD_10549 replaced by ADD_11602

//BasicMUL48_660 replaced by BasicMUL48_967

//BasicMUL48_661 replaced by BasicMUL48_958

//BasicMUL48_662 replaced by BasicMUL48_967

//ADD_10554 replaced by ADD_11595

//ADD_10553 replaced by ADD_11602

//ADD_10552 replaced by ADD_11602

//ADD_10557 replaced by ADD_11592

//ADD_10556 replaced by ADD_11602

//ADD_10555 replaced by ADD_11602

//ADD_10560 replaced by ADD_11592

//ADD_10559 replaced by ADD_11602

//ADD_10558 replaced by ADD_11602

//ADD_10563 replaced by ADD_11595

//ADD_10562 replaced by ADD_11602

//ADD_10561 replaced by ADD_11602

//BasicMUL48_663 replaced by BasicMUL48_970

//BasicMUL48_664 replaced by BasicMUL48_967

//BasicMUL48_665 replaced by BasicMUL48_970

//ADD_10566 replaced by ADD_11602

//ADD_10565 replaced by ADD_11602

//ADD_10564 replaced by ADD_11602

//ADD_10569 replaced by ADD_11601

//ADD_10568 replaced by ADD_11602

//ADD_10567 replaced by ADD_11602

//ADD_10571 replaced by ADD_11602

//ADD_10570 replaced by ADD_11602

//BasicMUL48_666 replaced by BasicMUL48_971

//BasicMUL48_667 replaced by BasicMUL48_970

//BasicMUL48_668 replaced by BasicMUL48_971

//ADD_10574 replaced by ADD_11595

//ADD_10573 replaced by ADD_11602

//ADD_10572 replaced by ADD_11602

//ADD_10577 replaced by ADD_11592

//ADD_10576 replaced by ADD_11602

//ADD_10575 replaced by ADD_11602

//ADD_10580 replaced by ADD_11592

//ADD_10579 replaced by ADD_11602

//ADD_10578 replaced by ADD_11602

//ADD_10583 replaced by ADD_11595

//ADD_10582 replaced by ADD_11602

//ADD_10581 replaced by ADD_11602

//BasicMUL48_669 replaced by BasicMUL48_970

//BasicMUL48_670 replaced by BasicMUL48_967

//BasicMUL48_671 replaced by BasicMUL48_970

//ADD_10586 replaced by ADD_11602

//ADD_10585 replaced by ADD_11602

//ADD_10584 replaced by ADD_11602

//ADD_10589 replaced by ADD_11601

//ADD_10588 replaced by ADD_11602

//ADD_10587 replaced by ADD_11602

//ADD_10591 replaced by ADD_11602

//ADD_10590 replaced by ADD_11602

//BasicMUL48_672 replaced by BasicMUL48_971

//BasicMUL48_673 replaced by BasicMUL48_970

//BasicMUL48_674 replaced by BasicMUL48_971

//ADD_10594 replaced by ADD_11602

//ADD_10593 replaced by ADD_11602

//ADD_10592 replaced by ADD_11602

//ADD_10597 replaced by ADD_11601

//ADD_10596 replaced by ADD_11602

//ADD_10595 replaced by ADD_11602

//ADD_10599 replaced by ADD_11602

//ADD_10598 replaced by ADD_11602

//BasicMUL48_675 replaced by BasicMUL48_971

//BasicMUL48_676 replaced by BasicMUL48_970

//BasicMUL48_677 replaced by BasicMUL48_971

//ADD_10602 replaced by ADD_11595

//ADD_10601 replaced by ADD_11602

//ADD_10600 replaced by ADD_11602

//ADD_10605 replaced by ADD_11592

//ADD_10604 replaced by ADD_11602

//ADD_10603 replaced by ADD_11602

//ADD_10608 replaced by ADD_11592

//ADD_10607 replaced by ADD_11602

//ADD_10606 replaced by ADD_11602

//ADD_10611 replaced by ADD_11595

//ADD_10610 replaced by ADD_11602

//ADD_10609 replaced by ADD_11602

//BasicMUL48_678 replaced by BasicMUL48_970

//BasicMUL48_679 replaced by BasicMUL48_967

//BasicMUL48_680 replaced by BasicMUL48_970

//ADD_10614 replaced by ADD_11602

//ADD_10613 replaced by ADD_11602

//ADD_10612 replaced by ADD_11602

//ADD_10617 replaced by ADD_11601

//ADD_10616 replaced by ADD_11602

//ADD_10615 replaced by ADD_11602

//ADD_10619 replaced by ADD_11602

//ADD_10618 replaced by ADD_11602

//BasicMUL48_681 replaced by BasicMUL48_971

//BasicMUL48_682 replaced by BasicMUL48_970

//BasicMUL48_683 replaced by BasicMUL48_971

//ADD_10622 replaced by ADD_11595

//ADD_10621 replaced by ADD_11602

//ADD_10620 replaced by ADD_11602

//ADD_10625 replaced by ADD_11592

//ADD_10624 replaced by ADD_11602

//ADD_10623 replaced by ADD_11602

//ADD_10628 replaced by ADD_11592

//ADD_10627 replaced by ADD_11602

//ADD_10626 replaced by ADD_11602

//ADD_10631 replaced by ADD_11595

//ADD_10630 replaced by ADD_11602

//ADD_10629 replaced by ADD_11602

//BasicMUL48_684 replaced by BasicMUL48_970

//BasicMUL48_685 replaced by BasicMUL48_967

//BasicMUL48_686 replaced by BasicMUL48_970

//ADD_10634 replaced by ADD_11563

//ADD_10633 replaced by ADD_11602

//ADD_10632 replaced by ADD_11602

//ADD_10637 replaced by ADD_11560

//ADD_10636 replaced by ADD_11602

//ADD_10635 replaced by ADD_11602

//ADD_10640 replaced by ADD_11560

//ADD_10639 replaced by ADD_11602

//ADD_10638 replaced by ADD_11602

//ADD_10643 replaced by ADD_11563

//ADD_10642 replaced by ADD_11602

//ADD_10641 replaced by ADD_11602

//BasicMUL48_687 replaced by BasicMUL48_967

//BasicMUL48_688 replaced by BasicMUL48_958

//BasicMUL48_689 replaced by BasicMUL48_967

//ADD_10646 replaced by ADD_11595

//ADD_10645 replaced by ADD_11602

//ADD_10644 replaced by ADD_11602

//ADD_10649 replaced by ADD_11592

//ADD_10648 replaced by ADD_11602

//ADD_10647 replaced by ADD_11602

//ADD_10652 replaced by ADD_11592

//ADD_10651 replaced by ADD_11602

//ADD_10650 replaced by ADD_11602

//ADD_10655 replaced by ADD_11595

//ADD_10654 replaced by ADD_11602

//ADD_10653 replaced by ADD_11602

//BasicMUL48_690 replaced by BasicMUL48_970

//BasicMUL48_691 replaced by BasicMUL48_967

//BasicMUL48_692 replaced by BasicMUL48_970

//ADD_10658 replaced by ADD_11602

//ADD_10657 replaced by ADD_11602

//ADD_10656 replaced by ADD_11602

//ADD_10661 replaced by ADD_11601

//ADD_10660 replaced by ADD_11602

//ADD_10659 replaced by ADD_11602

//ADD_10663 replaced by ADD_11602

//ADD_10662 replaced by ADD_11602

//BasicMUL48_693 replaced by BasicMUL48_971

//BasicMUL48_694 replaced by BasicMUL48_970

//BasicMUL48_695 replaced by BasicMUL48_971

//ADD_10666 replaced by ADD_11595

//ADD_10665 replaced by ADD_11602

//ADD_10664 replaced by ADD_11602

//ADD_10669 replaced by ADD_11592

//ADD_10668 replaced by ADD_11602

//ADD_10667 replaced by ADD_11602

//ADD_10672 replaced by ADD_11592

//ADD_10671 replaced by ADD_11602

//ADD_10670 replaced by ADD_11602

//ADD_10675 replaced by ADD_11595

//ADD_10674 replaced by ADD_11602

//ADD_10673 replaced by ADD_11602

//BasicMUL48_696 replaced by BasicMUL48_970

//BasicMUL48_697 replaced by BasicMUL48_967

//BasicMUL48_698 replaced by BasicMUL48_970

//ADD_10678 replaced by ADD_11602

//ADD_10677 replaced by ADD_11602

//ADD_10676 replaced by ADD_11602

//ADD_10681 replaced by ADD_11601

//ADD_10680 replaced by ADD_11602

//ADD_10679 replaced by ADD_11602

//ADD_10683 replaced by ADD_11602

//ADD_10682 replaced by ADD_11602

//BasicMUL48_699 replaced by BasicMUL48_971

//BasicMUL48_700 replaced by BasicMUL48_970

//BasicMUL48_701 replaced by BasicMUL48_971

//ADD_10686 replaced by ADD_11602

//ADD_10685 replaced by ADD_11602

//ADD_10684 replaced by ADD_11602

//ADD_10689 replaced by ADD_11601

//ADD_10688 replaced by ADD_11602

//ADD_10687 replaced by ADD_11602

//ADD_10691 replaced by ADD_11602

//ADD_10690 replaced by ADD_11602

//BasicMUL48_702 replaced by BasicMUL48_971

//BasicMUL48_703 replaced by BasicMUL48_970

//BasicMUL48_704 replaced by BasicMUL48_971

//ADD_10694 replaced by ADD_11595

//ADD_10693 replaced by ADD_11602

//ADD_10692 replaced by ADD_11602

//ADD_10697 replaced by ADD_11592

//ADD_10696 replaced by ADD_11602

//ADD_10695 replaced by ADD_11602

//ADD_10700 replaced by ADD_11592

//ADD_10699 replaced by ADD_11602

//ADD_10698 replaced by ADD_11602

//ADD_10703 replaced by ADD_11595

//ADD_10702 replaced by ADD_11602

//ADD_10701 replaced by ADD_11602

//BasicMUL48_705 replaced by BasicMUL48_970

//BasicMUL48_706 replaced by BasicMUL48_967

//BasicMUL48_707 replaced by BasicMUL48_970

//ADD_10706 replaced by ADD_11602

//ADD_10705 replaced by ADD_11602

//ADD_10704 replaced by ADD_11602

//ADD_10709 replaced by ADD_11601

//ADD_10708 replaced by ADD_11602

//ADD_10707 replaced by ADD_11602

//ADD_10711 replaced by ADD_11602

//ADD_10710 replaced by ADD_11602

//BasicMUL48_708 replaced by BasicMUL48_971

//BasicMUL48_709 replaced by BasicMUL48_970

//BasicMUL48_710 replaced by BasicMUL48_971

//ADD_10714 replaced by ADD_11595

//ADD_10713 replaced by ADD_11602

//ADD_10712 replaced by ADD_11602

//ADD_10717 replaced by ADD_11592

//ADD_10716 replaced by ADD_11602

//ADD_10715 replaced by ADD_11602

//ADD_10720 replaced by ADD_11592

//ADD_10719 replaced by ADD_11602

//ADD_10718 replaced by ADD_11602

//ADD_10723 replaced by ADD_11595

//ADD_10722 replaced by ADD_11602

//ADD_10721 replaced by ADD_11602

//BasicMUL48_711 replaced by BasicMUL48_970

//BasicMUL48_712 replaced by BasicMUL48_967

//BasicMUL48_713 replaced by BasicMUL48_970

//ADD_10726 replaced by ADD_11563

//ADD_10725 replaced by ADD_11602

//ADD_10724 replaced by ADD_11602

//ADD_10729 replaced by ADD_11560

//ADD_10728 replaced by ADD_11602

//ADD_10727 replaced by ADD_11602

//ADD_10732 replaced by ADD_11560

//ADD_10731 replaced by ADD_11602

//ADD_10730 replaced by ADD_11602

//ADD_10735 replaced by ADD_11563

//ADD_10734 replaced by ADD_11602

//ADD_10733 replaced by ADD_11602

//BasicMUL48_714 replaced by BasicMUL48_967

//BasicMUL48_715 replaced by BasicMUL48_958

//BasicMUL48_716 replaced by BasicMUL48_967

//ADD_10738 replaced by ADD_11595

//ADD_10737 replaced by ADD_11602

//ADD_10736 replaced by ADD_11602

//ADD_10741 replaced by ADD_11592

//ADD_10740 replaced by ADD_11602

//ADD_10739 replaced by ADD_11602

//ADD_10744 replaced by ADD_11592

//ADD_10743 replaced by ADD_11602

//ADD_10742 replaced by ADD_11602

//ADD_10747 replaced by ADD_11595

//ADD_10746 replaced by ADD_11602

//ADD_10745 replaced by ADD_11602

//BasicMUL48_717 replaced by BasicMUL48_970

//BasicMUL48_718 replaced by BasicMUL48_967

//BasicMUL48_719 replaced by BasicMUL48_970

//ADD_10750 replaced by ADD_11602

//ADD_10749 replaced by ADD_11602

//ADD_10748 replaced by ADD_11602

//ADD_10753 replaced by ADD_11601

//ADD_10752 replaced by ADD_11602

//ADD_10751 replaced by ADD_11602

//ADD_10755 replaced by ADD_11602

//ADD_10754 replaced by ADD_11602

//BasicMUL48_720 replaced by BasicMUL48_971

//BasicMUL48_721 replaced by BasicMUL48_970

//BasicMUL48_722 replaced by BasicMUL48_971

//ADD_10758 replaced by ADD_11595

//ADD_10757 replaced by ADD_11602

//ADD_10756 replaced by ADD_11602

//ADD_10761 replaced by ADD_11592

//ADD_10760 replaced by ADD_11602

//ADD_10759 replaced by ADD_11602

//ADD_10764 replaced by ADD_11592

//ADD_10763 replaced by ADD_11602

//ADD_10762 replaced by ADD_11602

//ADD_10767 replaced by ADD_11595

//ADD_10766 replaced by ADD_11602

//ADD_10765 replaced by ADD_11602

//BasicMUL48_723 replaced by BasicMUL48_970

//BasicMUL48_724 replaced by BasicMUL48_967

//BasicMUL48_725 replaced by BasicMUL48_970

//ADD_10770 replaced by ADD_11602

//ADD_10769 replaced by ADD_11602

//ADD_10768 replaced by ADD_11602

//ADD_10773 replaced by ADD_11601

//ADD_10772 replaced by ADD_11602

//ADD_10771 replaced by ADD_11602

//ADD_10775 replaced by ADD_11602

//ADD_10774 replaced by ADD_11602

//BasicMUL48_726 replaced by BasicMUL48_971

//BasicMUL48_727 replaced by BasicMUL48_970

//BasicMUL48_728 replaced by BasicMUL48_971

//ADD_10778 replaced by ADD_11602

//ADD_10777 replaced by ADD_11602

//ADD_10776 replaced by ADD_11602

//ADD_10781 replaced by ADD_11601

//ADD_10780 replaced by ADD_11602

//ADD_10779 replaced by ADD_11602

//ADD_10783 replaced by ADD_11602

//ADD_10782 replaced by ADD_11602

//BasicMUL48_729 replaced by BasicMUL48_971

//BasicMUL48_730 replaced by BasicMUL48_970

//BasicMUL48_731 replaced by BasicMUL48_971

//ADD_10786 replaced by ADD_11595

//ADD_10785 replaced by ADD_11602

//ADD_10784 replaced by ADD_11602

//ADD_10789 replaced by ADD_11592

//ADD_10788 replaced by ADD_11602

//ADD_10787 replaced by ADD_11602

//ADD_10792 replaced by ADD_11592

//ADD_10791 replaced by ADD_11602

//ADD_10790 replaced by ADD_11602

//ADD_10795 replaced by ADD_11595

//ADD_10794 replaced by ADD_11602

//ADD_10793 replaced by ADD_11602

//BasicMUL48_732 replaced by BasicMUL48_970

//BasicMUL48_733 replaced by BasicMUL48_967

//BasicMUL48_734 replaced by BasicMUL48_970

//ADD_10798 replaced by ADD_11602

//ADD_10797 replaced by ADD_11602

//ADD_10796 replaced by ADD_11602

//ADD_10801 replaced by ADD_11601

//ADD_10800 replaced by ADD_11602

//ADD_10799 replaced by ADD_11602

//ADD_10803 replaced by ADD_11602

//ADD_10802 replaced by ADD_11602

//BasicMUL48_735 replaced by BasicMUL48_971

//BasicMUL48_736 replaced by BasicMUL48_970

//BasicMUL48_737 replaced by BasicMUL48_971

//ADD_10806 replaced by ADD_11595

//ADD_10805 replaced by ADD_11602

//ADD_10804 replaced by ADD_11602

//ADD_10809 replaced by ADD_11592

//ADD_10808 replaced by ADD_11602

//ADD_10807 replaced by ADD_11602

//ADD_10812 replaced by ADD_11592

//ADD_10811 replaced by ADD_11602

//ADD_10810 replaced by ADD_11602

//ADD_10815 replaced by ADD_11595

//ADD_10814 replaced by ADD_11602

//ADD_10813 replaced by ADD_11602

//BasicMUL48_738 replaced by BasicMUL48_970

//BasicMUL48_739 replaced by BasicMUL48_967

//BasicMUL48_740 replaced by BasicMUL48_970

//ADD_10818 replaced by ADD_11563

//ADD_10817 replaced by ADD_11602

//ADD_10816 replaced by ADD_11602

//ADD_10821 replaced by ADD_11560

//ADD_10820 replaced by ADD_11602

//ADD_10819 replaced by ADD_11602

//ADD_10824 replaced by ADD_11560

//ADD_10823 replaced by ADD_11602

//ADD_10822 replaced by ADD_11602

//ADD_10827 replaced by ADD_11563

//ADD_10826 replaced by ADD_11602

//ADD_10825 replaced by ADD_11602

//BasicMUL48_741 replaced by BasicMUL48_967

//BasicMUL48_742 replaced by BasicMUL48_958

//BasicMUL48_743 replaced by BasicMUL48_967

//ADD_10830 replaced by ADD_11595

//ADD_10829 replaced by ADD_11602

//ADD_10828 replaced by ADD_11602

//ADD_10833 replaced by ADD_11592

//ADD_10832 replaced by ADD_11602

//ADD_10831 replaced by ADD_11602

//ADD_10836 replaced by ADD_11592

//ADD_10835 replaced by ADD_11602

//ADD_10834 replaced by ADD_11602

//ADD_10839 replaced by ADD_11595

//ADD_10838 replaced by ADD_11602

//ADD_10837 replaced by ADD_11602

//BasicMUL48_744 replaced by BasicMUL48_970

//BasicMUL48_745 replaced by BasicMUL48_967

//BasicMUL48_746 replaced by BasicMUL48_970

//ADD_10842 replaced by ADD_11602

//ADD_10841 replaced by ADD_11602

//ADD_10840 replaced by ADD_11602

//ADD_10845 replaced by ADD_11601

//ADD_10844 replaced by ADD_11602

//ADD_10843 replaced by ADD_11602

//ADD_10847 replaced by ADD_11602

//ADD_10846 replaced by ADD_11602

//BasicMUL48_747 replaced by BasicMUL48_971

//BasicMUL48_748 replaced by BasicMUL48_970

//BasicMUL48_749 replaced by BasicMUL48_971

//ADD_10850 replaced by ADD_11595

//ADD_10849 replaced by ADD_11602

//ADD_10848 replaced by ADD_11602

//ADD_10853 replaced by ADD_11592

//ADD_10852 replaced by ADD_11602

//ADD_10851 replaced by ADD_11602

//ADD_10856 replaced by ADD_11592

//ADD_10855 replaced by ADD_11602

//ADD_10854 replaced by ADD_11602

//ADD_10859 replaced by ADD_11595

//ADD_10858 replaced by ADD_11602

//ADD_10857 replaced by ADD_11602

//BasicMUL48_750 replaced by BasicMUL48_970

//BasicMUL48_751 replaced by BasicMUL48_967

//BasicMUL48_752 replaced by BasicMUL48_970

//ADD_10862 replaced by ADD_11602

//ADD_10861 replaced by ADD_11602

//ADD_10860 replaced by ADD_11602

//ADD_10865 replaced by ADD_11601

//ADD_10864 replaced by ADD_11602

//ADD_10863 replaced by ADD_11602

//ADD_10867 replaced by ADD_11602

//ADD_10866 replaced by ADD_11602

//BasicMUL48_753 replaced by BasicMUL48_971

//BasicMUL48_754 replaced by BasicMUL48_970

//BasicMUL48_755 replaced by BasicMUL48_971

//ADD_10870 replaced by ADD_11602

//ADD_10869 replaced by ADD_11602

//ADD_10868 replaced by ADD_11602

//ADD_10873 replaced by ADD_11601

//ADD_10872 replaced by ADD_11602

//ADD_10871 replaced by ADD_11602

//ADD_10875 replaced by ADD_11602

//ADD_10874 replaced by ADD_11602

//BasicMUL48_756 replaced by BasicMUL48_971

//BasicMUL48_757 replaced by BasicMUL48_970

//BasicMUL48_758 replaced by BasicMUL48_971

//ADD_10878 replaced by ADD_11595

//ADD_10877 replaced by ADD_11602

//ADD_10876 replaced by ADD_11602

//ADD_10881 replaced by ADD_11592

//ADD_10880 replaced by ADD_11602

//ADD_10879 replaced by ADD_11602

//ADD_10884 replaced by ADD_11592

//ADD_10883 replaced by ADD_11602

//ADD_10882 replaced by ADD_11602

//ADD_10887 replaced by ADD_11595

//ADD_10886 replaced by ADD_11602

//ADD_10885 replaced by ADD_11602

//BasicMUL48_759 replaced by BasicMUL48_970

//BasicMUL48_760 replaced by BasicMUL48_967

//BasicMUL48_761 replaced by BasicMUL48_970

//ADD_10890 replaced by ADD_11602

//ADD_10889 replaced by ADD_11602

//ADD_10888 replaced by ADD_11602

//ADD_10893 replaced by ADD_11601

//ADD_10892 replaced by ADD_11602

//ADD_10891 replaced by ADD_11602

//ADD_10895 replaced by ADD_11602

//ADD_10894 replaced by ADD_11602

//BasicMUL48_762 replaced by BasicMUL48_971

//BasicMUL48_763 replaced by BasicMUL48_970

//BasicMUL48_764 replaced by BasicMUL48_971

//ADD_10898 replaced by ADD_11595

//ADD_10897 replaced by ADD_11602

//ADD_10896 replaced by ADD_11602

//ADD_10901 replaced by ADD_11592

//ADD_10900 replaced by ADD_11602

//ADD_10899 replaced by ADD_11602

//ADD_10904 replaced by ADD_11592

//ADD_10903 replaced by ADD_11602

//ADD_10902 replaced by ADD_11602

//ADD_10907 replaced by ADD_11595

//ADD_10906 replaced by ADD_11602

//ADD_10905 replaced by ADD_11602

//BasicMUL48_765 replaced by BasicMUL48_970

//BasicMUL48_766 replaced by BasicMUL48_967

//BasicMUL48_767 replaced by BasicMUL48_970

//ADD_10910 replaced by ADD_11563

//ADD_10909 replaced by ADD_11602

//ADD_10908 replaced by ADD_11602

//ADD_10913 replaced by ADD_11560

//ADD_10912 replaced by ADD_11602

//ADD_10911 replaced by ADD_11602

//ADD_10916 replaced by ADD_11560

//ADD_10915 replaced by ADD_11602

//ADD_10914 replaced by ADD_11602

//ADD_10919 replaced by ADD_11563

//ADD_10918 replaced by ADD_11602

//ADD_10917 replaced by ADD_11602

//BasicMUL48_768 replaced by BasicMUL48_967

//BasicMUL48_769 replaced by BasicMUL48_958

//BasicMUL48_770 replaced by BasicMUL48_967

//ADD_10922 replaced by ADD_11595

//ADD_10921 replaced by ADD_11602

//ADD_10920 replaced by ADD_11602

//ADD_10925 replaced by ADD_11592

//ADD_10924 replaced by ADD_11602

//ADD_10923 replaced by ADD_11602

//ADD_10928 replaced by ADD_11592

//ADD_10927 replaced by ADD_11602

//ADD_10926 replaced by ADD_11602

//ADD_10931 replaced by ADD_11595

//ADD_10930 replaced by ADD_11602

//ADD_10929 replaced by ADD_11602

//BasicMUL48_771 replaced by BasicMUL48_970

//BasicMUL48_772 replaced by BasicMUL48_967

//BasicMUL48_773 replaced by BasicMUL48_970

//ADD_10934 replaced by ADD_11602

//ADD_10933 replaced by ADD_11602

//ADD_10932 replaced by ADD_11602

//ADD_10937 replaced by ADD_11601

//ADD_10936 replaced by ADD_11602

//ADD_10935 replaced by ADD_11602

//ADD_10939 replaced by ADD_11602

//ADD_10938 replaced by ADD_11602

//BasicMUL48_774 replaced by BasicMUL48_971

//BasicMUL48_775 replaced by BasicMUL48_970

//BasicMUL48_776 replaced by BasicMUL48_971

//ADD_10942 replaced by ADD_11595

//ADD_10941 replaced by ADD_11602

//ADD_10940 replaced by ADD_11602

//ADD_10945 replaced by ADD_11592

//ADD_10944 replaced by ADD_11602

//ADD_10943 replaced by ADD_11602

//ADD_10948 replaced by ADD_11592

//ADD_10947 replaced by ADD_11602

//ADD_10946 replaced by ADD_11602

//ADD_10951 replaced by ADD_11595

//ADD_10950 replaced by ADD_11602

//ADD_10949 replaced by ADD_11602

//BasicMUL48_777 replaced by BasicMUL48_970

//BasicMUL48_778 replaced by BasicMUL48_967

//BasicMUL48_779 replaced by BasicMUL48_970

//ADD_10954 replaced by ADD_11602

//ADD_10953 replaced by ADD_11602

//ADD_10952 replaced by ADD_11602

//ADD_10957 replaced by ADD_11601

//ADD_10956 replaced by ADD_11602

//ADD_10955 replaced by ADD_11602

//ADD_10959 replaced by ADD_11602

//ADD_10958 replaced by ADD_11602

//BasicMUL48_780 replaced by BasicMUL48_971

//BasicMUL48_781 replaced by BasicMUL48_970

//BasicMUL48_782 replaced by BasicMUL48_971

//ADD_10962 replaced by ADD_11602

//ADD_10961 replaced by ADD_11602

//ADD_10960 replaced by ADD_11602

//ADD_10965 replaced by ADD_11601

//ADD_10964 replaced by ADD_11602

//ADD_10963 replaced by ADD_11602

//ADD_10967 replaced by ADD_11602

//ADD_10966 replaced by ADD_11602

//BasicMUL48_783 replaced by BasicMUL48_971

//BasicMUL48_784 replaced by BasicMUL48_970

//BasicMUL48_785 replaced by BasicMUL48_971

//ADD_10970 replaced by ADD_11595

//ADD_10969 replaced by ADD_11602

//ADD_10968 replaced by ADD_11602

//ADD_10973 replaced by ADD_11592

//ADD_10972 replaced by ADD_11602

//ADD_10971 replaced by ADD_11602

//ADD_10976 replaced by ADD_11592

//ADD_10975 replaced by ADD_11602

//ADD_10974 replaced by ADD_11602

//ADD_10979 replaced by ADD_11595

//ADD_10978 replaced by ADD_11602

//ADD_10977 replaced by ADD_11602

//BasicMUL48_786 replaced by BasicMUL48_970

//BasicMUL48_787 replaced by BasicMUL48_967

//BasicMUL48_788 replaced by BasicMUL48_970

//ADD_10982 replaced by ADD_11602

//ADD_10981 replaced by ADD_11602

//ADD_10980 replaced by ADD_11602

//ADD_10985 replaced by ADD_11601

//ADD_10984 replaced by ADD_11602

//ADD_10983 replaced by ADD_11602

//ADD_10987 replaced by ADD_11602

//ADD_10986 replaced by ADD_11602

//BasicMUL48_789 replaced by BasicMUL48_971

//BasicMUL48_790 replaced by BasicMUL48_970

//BasicMUL48_791 replaced by BasicMUL48_971

//ADD_10990 replaced by ADD_11595

//ADD_10989 replaced by ADD_11602

//ADD_10988 replaced by ADD_11602

//ADD_10993 replaced by ADD_11592

//ADD_10992 replaced by ADD_11602

//ADD_10991 replaced by ADD_11602

//ADD_10996 replaced by ADD_11592

//ADD_10995 replaced by ADD_11602

//ADD_10994 replaced by ADD_11602

//ADD_10999 replaced by ADD_11595

//ADD_10998 replaced by ADD_11602

//ADD_10997 replaced by ADD_11602

//BasicMUL48_792 replaced by BasicMUL48_970

//BasicMUL48_793 replaced by BasicMUL48_967

//BasicMUL48_794 replaced by BasicMUL48_970

//ADD_11002 replaced by ADD_11563

//ADD_11001 replaced by ADD_11602

//ADD_11000 replaced by ADD_11602

//ADD_11005 replaced by ADD_11560

//ADD_11004 replaced by ADD_11602

//ADD_11003 replaced by ADD_11602

//ADD_11008 replaced by ADD_11560

//ADD_11007 replaced by ADD_11602

//ADD_11006 replaced by ADD_11602

//ADD_11011 replaced by ADD_11563

//ADD_11010 replaced by ADD_11602

//ADD_11009 replaced by ADD_11602

//BasicMUL48_795 replaced by BasicMUL48_967

//BasicMUL48_796 replaced by BasicMUL48_958

//BasicMUL48_797 replaced by BasicMUL48_967

//ADD_11014 replaced by ADD_11595

//ADD_11013 replaced by ADD_11602

//ADD_11012 replaced by ADD_11602

//ADD_11017 replaced by ADD_11592

//ADD_11016 replaced by ADD_11602

//ADD_11015 replaced by ADD_11602

//ADD_11020 replaced by ADD_11592

//ADD_11019 replaced by ADD_11602

//ADD_11018 replaced by ADD_11602

//ADD_11023 replaced by ADD_11595

//ADD_11022 replaced by ADD_11602

//ADD_11021 replaced by ADD_11602

//BasicMUL48_798 replaced by BasicMUL48_970

//BasicMUL48_799 replaced by BasicMUL48_967

//BasicMUL48_800 replaced by BasicMUL48_970

//ADD_11026 replaced by ADD_11602

//ADD_11025 replaced by ADD_11602

//ADD_11024 replaced by ADD_11602

//ADD_11029 replaced by ADD_11601

//ADD_11028 replaced by ADD_11602

//ADD_11027 replaced by ADD_11602

//ADD_11031 replaced by ADD_11602

//ADD_11030 replaced by ADD_11602

//BasicMUL48_801 replaced by BasicMUL48_971

//BasicMUL48_802 replaced by BasicMUL48_970

//BasicMUL48_803 replaced by BasicMUL48_971

//ADD_11034 replaced by ADD_11595

//ADD_11033 replaced by ADD_11602

//ADD_11032 replaced by ADD_11602

//ADD_11037 replaced by ADD_11592

//ADD_11036 replaced by ADD_11602

//ADD_11035 replaced by ADD_11602

//ADD_11040 replaced by ADD_11592

//ADD_11039 replaced by ADD_11602

//ADD_11038 replaced by ADD_11602

//ADD_11043 replaced by ADD_11595

//ADD_11042 replaced by ADD_11602

//ADD_11041 replaced by ADD_11602

//BasicMUL48_804 replaced by BasicMUL48_970

//BasicMUL48_805 replaced by BasicMUL48_967

//BasicMUL48_806 replaced by BasicMUL48_970

//ADD_11046 replaced by ADD_11602

//ADD_11045 replaced by ADD_11602

//ADD_11044 replaced by ADD_11602

//ADD_11049 replaced by ADD_11601

//ADD_11048 replaced by ADD_11602

//ADD_11047 replaced by ADD_11602

//ADD_11051 replaced by ADD_11602

//ADD_11050 replaced by ADD_11602

//BasicMUL48_807 replaced by BasicMUL48_971

//BasicMUL48_808 replaced by BasicMUL48_970

//BasicMUL48_809 replaced by BasicMUL48_971

//ADD_11054 replaced by ADD_11602

//ADD_11053 replaced by ADD_11602

//ADD_11052 replaced by ADD_11602

//ADD_11057 replaced by ADD_11601

//ADD_11056 replaced by ADD_11602

//ADD_11055 replaced by ADD_11602

//ADD_11059 replaced by ADD_11602

//ADD_11058 replaced by ADD_11602

//BasicMUL48_810 replaced by BasicMUL48_971

//BasicMUL48_811 replaced by BasicMUL48_970

//BasicMUL48_812 replaced by BasicMUL48_971

//ADD_11062 replaced by ADD_11595

//ADD_11061 replaced by ADD_11602

//ADD_11060 replaced by ADD_11602

//ADD_11065 replaced by ADD_11592

//ADD_11064 replaced by ADD_11602

//ADD_11063 replaced by ADD_11602

//ADD_11068 replaced by ADD_11592

//ADD_11067 replaced by ADD_11602

//ADD_11066 replaced by ADD_11602

//ADD_11071 replaced by ADD_11595

//ADD_11070 replaced by ADD_11602

//ADD_11069 replaced by ADD_11602

//BasicMUL48_813 replaced by BasicMUL48_970

//BasicMUL48_814 replaced by BasicMUL48_967

//BasicMUL48_815 replaced by BasicMUL48_970

//ADD_11074 replaced by ADD_11602

//ADD_11073 replaced by ADD_11602

//ADD_11072 replaced by ADD_11602

//ADD_11077 replaced by ADD_11601

//ADD_11076 replaced by ADD_11602

//ADD_11075 replaced by ADD_11602

//ADD_11079 replaced by ADD_11602

//ADD_11078 replaced by ADD_11602

//BasicMUL48_816 replaced by BasicMUL48_971

//BasicMUL48_817 replaced by BasicMUL48_970

//BasicMUL48_818 replaced by BasicMUL48_971

//ADD_11082 replaced by ADD_11595

//ADD_11081 replaced by ADD_11602

//ADD_11080 replaced by ADD_11602

//ADD_11085 replaced by ADD_11592

//ADD_11084 replaced by ADD_11602

//ADD_11083 replaced by ADD_11602

//ADD_11088 replaced by ADD_11592

//ADD_11087 replaced by ADD_11602

//ADD_11086 replaced by ADD_11602

//ADD_11091 replaced by ADD_11595

//ADD_11090 replaced by ADD_11602

//ADD_11089 replaced by ADD_11602

//BasicMUL48_819 replaced by BasicMUL48_970

//BasicMUL48_820 replaced by BasicMUL48_967

//BasicMUL48_821 replaced by BasicMUL48_970

//ADD_11094 replaced by ADD_11563

//ADD_11093 replaced by ADD_11602

//ADD_11092 replaced by ADD_11602

//ADD_11097 replaced by ADD_11560

//ADD_11096 replaced by ADD_11602

//ADD_11095 replaced by ADD_11602

//ADD_11100 replaced by ADD_11560

//ADD_11099 replaced by ADD_11602

//ADD_11098 replaced by ADD_11602

//ADD_11103 replaced by ADD_11563

//ADD_11102 replaced by ADD_11602

//ADD_11101 replaced by ADD_11602

//BasicMUL48_822 replaced by BasicMUL48_967

//BasicMUL48_823 replaced by BasicMUL48_958

//BasicMUL48_824 replaced by BasicMUL48_967

//ADD_11106 replaced by ADD_11595

//ADD_11105 replaced by ADD_11602

//ADD_11104 replaced by ADD_11602

//ADD_11109 replaced by ADD_11592

//ADD_11108 replaced by ADD_11602

//ADD_11107 replaced by ADD_11602

//ADD_11112 replaced by ADD_11592

//ADD_11111 replaced by ADD_11602

//ADD_11110 replaced by ADD_11602

//ADD_11115 replaced by ADD_11595

//ADD_11114 replaced by ADD_11602

//ADD_11113 replaced by ADD_11602

//BasicMUL48_825 replaced by BasicMUL48_970

//BasicMUL48_826 replaced by BasicMUL48_967

//BasicMUL48_827 replaced by BasicMUL48_970

//ADD_11118 replaced by ADD_11602

//ADD_11117 replaced by ADD_11602

//ADD_11116 replaced by ADD_11602

//ADD_11121 replaced by ADD_11601

//ADD_11120 replaced by ADD_11602

//ADD_11119 replaced by ADD_11602

//ADD_11123 replaced by ADD_11602

//ADD_11122 replaced by ADD_11602

//BasicMUL48_828 replaced by BasicMUL48_971

//BasicMUL48_829 replaced by BasicMUL48_970

//BasicMUL48_830 replaced by BasicMUL48_971

//ADD_11126 replaced by ADD_11595

//ADD_11125 replaced by ADD_11602

//ADD_11124 replaced by ADD_11602

//ADD_11129 replaced by ADD_11592

//ADD_11128 replaced by ADD_11602

//ADD_11127 replaced by ADD_11602

//ADD_11132 replaced by ADD_11592

//ADD_11131 replaced by ADD_11602

//ADD_11130 replaced by ADD_11602

//ADD_11135 replaced by ADD_11595

//ADD_11134 replaced by ADD_11602

//ADD_11133 replaced by ADD_11602

//BasicMUL48_831 replaced by BasicMUL48_970

//BasicMUL48_832 replaced by BasicMUL48_967

//BasicMUL48_833 replaced by BasicMUL48_970

//ADD_11138 replaced by ADD_11602

//ADD_11137 replaced by ADD_11602

//ADD_11136 replaced by ADD_11602

//ADD_11141 replaced by ADD_11601

//ADD_11140 replaced by ADD_11602

//ADD_11139 replaced by ADD_11602

//ADD_11143 replaced by ADD_11602

//ADD_11142 replaced by ADD_11602

//BasicMUL48_834 replaced by BasicMUL48_971

//BasicMUL48_835 replaced by BasicMUL48_970

//BasicMUL48_836 replaced by BasicMUL48_971

//ADD_11146 replaced by ADD_11602

//ADD_11145 replaced by ADD_11602

//ADD_11144 replaced by ADD_11602

//ADD_11149 replaced by ADD_11601

//ADD_11148 replaced by ADD_11602

//ADD_11147 replaced by ADD_11602

//ADD_11151 replaced by ADD_11602

//ADD_11150 replaced by ADD_11602

//BasicMUL48_837 replaced by BasicMUL48_971

//BasicMUL48_838 replaced by BasicMUL48_970

//BasicMUL48_839 replaced by BasicMUL48_971

//ADD_11154 replaced by ADD_11595

//ADD_11153 replaced by ADD_11602

//ADD_11152 replaced by ADD_11602

//ADD_11157 replaced by ADD_11592

//ADD_11156 replaced by ADD_11602

//ADD_11155 replaced by ADD_11602

//ADD_11160 replaced by ADD_11592

//ADD_11159 replaced by ADD_11602

//ADD_11158 replaced by ADD_11602

//ADD_11163 replaced by ADD_11595

//ADD_11162 replaced by ADD_11602

//ADD_11161 replaced by ADD_11602

//BasicMUL48_840 replaced by BasicMUL48_970

//BasicMUL48_841 replaced by BasicMUL48_967

//BasicMUL48_842 replaced by BasicMUL48_970

//ADD_11166 replaced by ADD_11602

//ADD_11165 replaced by ADD_11602

//ADD_11164 replaced by ADD_11602

//ADD_11169 replaced by ADD_11601

//ADD_11168 replaced by ADD_11602

//ADD_11167 replaced by ADD_11602

//ADD_11171 replaced by ADD_11602

//ADD_11170 replaced by ADD_11602

//BasicMUL48_843 replaced by BasicMUL48_971

//BasicMUL48_844 replaced by BasicMUL48_970

//BasicMUL48_845 replaced by BasicMUL48_971

//ADD_11174 replaced by ADD_11595

//ADD_11173 replaced by ADD_11602

//ADD_11172 replaced by ADD_11602

//ADD_11177 replaced by ADD_11592

//ADD_11176 replaced by ADD_11602

//ADD_11175 replaced by ADD_11602

//ADD_11180 replaced by ADD_11592

//ADD_11179 replaced by ADD_11602

//ADD_11178 replaced by ADD_11602

//ADD_11183 replaced by ADD_11595

//ADD_11182 replaced by ADD_11602

//ADD_11181 replaced by ADD_11602

//BasicMUL48_846 replaced by BasicMUL48_970

//BasicMUL48_847 replaced by BasicMUL48_967

//BasicMUL48_848 replaced by BasicMUL48_970

//ADD_11186 replaced by ADD_11563

//ADD_11185 replaced by ADD_11602

//ADD_11184 replaced by ADD_11602

//ADD_11189 replaced by ADD_11560

//ADD_11188 replaced by ADD_11602

//ADD_11187 replaced by ADD_11602

//ADD_11192 replaced by ADD_11560

//ADD_11191 replaced by ADD_11602

//ADD_11190 replaced by ADD_11602

//ADD_11195 replaced by ADD_11563

//ADD_11194 replaced by ADD_11602

//ADD_11193 replaced by ADD_11602

//BasicMUL48_849 replaced by BasicMUL48_967

//BasicMUL48_850 replaced by BasicMUL48_958

//BasicMUL48_851 replaced by BasicMUL48_967

//ADD_11198 replaced by ADD_11595

//ADD_11197 replaced by ADD_11602

//ADD_11196 replaced by ADD_11602

//ADD_11201 replaced by ADD_11592

//ADD_11200 replaced by ADD_11602

//ADD_11199 replaced by ADD_11602

//ADD_11204 replaced by ADD_11592

//ADD_11203 replaced by ADD_11602

//ADD_11202 replaced by ADD_11602

//ADD_11207 replaced by ADD_11595

//ADD_11206 replaced by ADD_11602

//ADD_11205 replaced by ADD_11602

//BasicMUL48_852 replaced by BasicMUL48_970

//BasicMUL48_853 replaced by BasicMUL48_967

//BasicMUL48_854 replaced by BasicMUL48_970

//ADD_11210 replaced by ADD_11602

//ADD_11209 replaced by ADD_11602

//ADD_11208 replaced by ADD_11602

//ADD_11213 replaced by ADD_11601

//ADD_11212 replaced by ADD_11602

//ADD_11211 replaced by ADD_11602

//ADD_11215 replaced by ADD_11602

//ADD_11214 replaced by ADD_11602

//BasicMUL48_855 replaced by BasicMUL48_971

//BasicMUL48_856 replaced by BasicMUL48_970

//BasicMUL48_857 replaced by BasicMUL48_971

//ADD_11218 replaced by ADD_11595

//ADD_11217 replaced by ADD_11602

//ADD_11216 replaced by ADD_11602

//ADD_11221 replaced by ADD_11592

//ADD_11220 replaced by ADD_11602

//ADD_11219 replaced by ADD_11602

//ADD_11224 replaced by ADD_11592

//ADD_11223 replaced by ADD_11602

//ADD_11222 replaced by ADD_11602

//ADD_11227 replaced by ADD_11595

//ADD_11226 replaced by ADD_11602

//ADD_11225 replaced by ADD_11602

//BasicMUL48_858 replaced by BasicMUL48_970

//BasicMUL48_859 replaced by BasicMUL48_967

//BasicMUL48_860 replaced by BasicMUL48_970

//ADD_11230 replaced by ADD_11602

//ADD_11229 replaced by ADD_11602

//ADD_11228 replaced by ADD_11602

//ADD_11233 replaced by ADD_11601

//ADD_11232 replaced by ADD_11602

//ADD_11231 replaced by ADD_11602

//ADD_11235 replaced by ADD_11602

//ADD_11234 replaced by ADD_11602

//BasicMUL48_861 replaced by BasicMUL48_971

//BasicMUL48_862 replaced by BasicMUL48_970

//BasicMUL48_863 replaced by BasicMUL48_971

//ADD_11238 replaced by ADD_11602

//ADD_11237 replaced by ADD_11602

//ADD_11236 replaced by ADD_11602

//ADD_11241 replaced by ADD_11601

//ADD_11240 replaced by ADD_11602

//ADD_11239 replaced by ADD_11602

//ADD_11243 replaced by ADD_11602

//ADD_11242 replaced by ADD_11602

//BasicMUL48_864 replaced by BasicMUL48_971

//BasicMUL48_865 replaced by BasicMUL48_970

//BasicMUL48_866 replaced by BasicMUL48_971

//ADD_11246 replaced by ADD_11595

//ADD_11245 replaced by ADD_11602

//ADD_11244 replaced by ADD_11602

//ADD_11249 replaced by ADD_11592

//ADD_11248 replaced by ADD_11602

//ADD_11247 replaced by ADD_11602

//ADD_11252 replaced by ADD_11592

//ADD_11251 replaced by ADD_11602

//ADD_11250 replaced by ADD_11602

//ADD_11255 replaced by ADD_11595

//ADD_11254 replaced by ADD_11602

//ADD_11253 replaced by ADD_11602

//BasicMUL48_867 replaced by BasicMUL48_970

//BasicMUL48_868 replaced by BasicMUL48_967

//BasicMUL48_869 replaced by BasicMUL48_970

//ADD_11258 replaced by ADD_11602

//ADD_11257 replaced by ADD_11602

//ADD_11256 replaced by ADD_11602

//ADD_11261 replaced by ADD_11601

//ADD_11260 replaced by ADD_11602

//ADD_11259 replaced by ADD_11602

//ADD_11263 replaced by ADD_11602

//ADD_11262 replaced by ADD_11602

//BasicMUL48_870 replaced by BasicMUL48_971

//BasicMUL48_871 replaced by BasicMUL48_970

//BasicMUL48_872 replaced by BasicMUL48_971

//ADD_11266 replaced by ADD_11595

//ADD_11265 replaced by ADD_11602

//ADD_11264 replaced by ADD_11602

//ADD_11269 replaced by ADD_11592

//ADD_11268 replaced by ADD_11602

//ADD_11267 replaced by ADD_11602

//ADD_11272 replaced by ADD_11592

//ADD_11271 replaced by ADD_11602

//ADD_11270 replaced by ADD_11602

//ADD_11275 replaced by ADD_11595

//ADD_11274 replaced by ADD_11602

//ADD_11273 replaced by ADD_11602

//BasicMUL48_873 replaced by BasicMUL48_970

//BasicMUL48_874 replaced by BasicMUL48_967

//BasicMUL48_875 replaced by BasicMUL48_970

//ADD_11278 replaced by ADD_11563

//ADD_11277 replaced by ADD_11602

//ADD_11276 replaced by ADD_11602

//ADD_11281 replaced by ADD_11560

//ADD_11280 replaced by ADD_11602

//ADD_11279 replaced by ADD_11602

//ADD_11284 replaced by ADD_11560

//ADD_11283 replaced by ADD_11602

//ADD_11282 replaced by ADD_11602

//ADD_11287 replaced by ADD_11563

//ADD_11286 replaced by ADD_11602

//ADD_11285 replaced by ADD_11602

//BasicMUL48_876 replaced by BasicMUL48_967

//BasicMUL48_877 replaced by BasicMUL48_958

//BasicMUL48_878 replaced by BasicMUL48_967

//ADD_11290 replaced by ADD_11595

//ADD_11289 replaced by ADD_11602

//ADD_11288 replaced by ADD_11602

//ADD_11293 replaced by ADD_11592

//ADD_11292 replaced by ADD_11602

//ADD_11291 replaced by ADD_11602

//ADD_11296 replaced by ADD_11592

//ADD_11295 replaced by ADD_11602

//ADD_11294 replaced by ADD_11602

//ADD_11299 replaced by ADD_11595

//ADD_11298 replaced by ADD_11602

//ADD_11297 replaced by ADD_11602

//BasicMUL48_879 replaced by BasicMUL48_970

//BasicMUL48_880 replaced by BasicMUL48_967

//BasicMUL48_881 replaced by BasicMUL48_970

//ADD_11302 replaced by ADD_11602

//ADD_11301 replaced by ADD_11602

//ADD_11300 replaced by ADD_11602

//ADD_11305 replaced by ADD_11601

//ADD_11304 replaced by ADD_11602

//ADD_11303 replaced by ADD_11602

//ADD_11307 replaced by ADD_11602

//ADD_11306 replaced by ADD_11602

//BasicMUL48_882 replaced by BasicMUL48_971

//BasicMUL48_883 replaced by BasicMUL48_970

//BasicMUL48_884 replaced by BasicMUL48_971

//ADD_11310 replaced by ADD_11595

//ADD_11309 replaced by ADD_11602

//ADD_11308 replaced by ADD_11602

//ADD_11313 replaced by ADD_11592

//ADD_11312 replaced by ADD_11602

//ADD_11311 replaced by ADD_11602

//ADD_11316 replaced by ADD_11592

//ADD_11315 replaced by ADD_11602

//ADD_11314 replaced by ADD_11602

//ADD_11319 replaced by ADD_11595

//ADD_11318 replaced by ADD_11602

//ADD_11317 replaced by ADD_11602

//BasicMUL48_885 replaced by BasicMUL48_970

//BasicMUL48_886 replaced by BasicMUL48_967

//BasicMUL48_887 replaced by BasicMUL48_970

//ADD_11322 replaced by ADD_11602

//ADD_11321 replaced by ADD_11602

//ADD_11320 replaced by ADD_11602

//ADD_11325 replaced by ADD_11601

//ADD_11324 replaced by ADD_11602

//ADD_11323 replaced by ADD_11602

//ADD_11327 replaced by ADD_11602

//ADD_11326 replaced by ADD_11602

//BasicMUL48_888 replaced by BasicMUL48_971

//BasicMUL48_889 replaced by BasicMUL48_970

//BasicMUL48_890 replaced by BasicMUL48_971

//ADD_11330 replaced by ADD_11602

//ADD_11329 replaced by ADD_11602

//ADD_11328 replaced by ADD_11602

//ADD_11333 replaced by ADD_11601

//ADD_11332 replaced by ADD_11602

//ADD_11331 replaced by ADD_11602

//ADD_11335 replaced by ADD_11602

//ADD_11334 replaced by ADD_11602

//BasicMUL48_891 replaced by BasicMUL48_971

//BasicMUL48_892 replaced by BasicMUL48_970

//BasicMUL48_893 replaced by BasicMUL48_971

//ADD_11338 replaced by ADD_11595

//ADD_11337 replaced by ADD_11602

//ADD_11336 replaced by ADD_11602

//ADD_11341 replaced by ADD_11592

//ADD_11340 replaced by ADD_11602

//ADD_11339 replaced by ADD_11602

//ADD_11344 replaced by ADD_11592

//ADD_11343 replaced by ADD_11602

//ADD_11342 replaced by ADD_11602

//ADD_11347 replaced by ADD_11595

//ADD_11346 replaced by ADD_11602

//ADD_11345 replaced by ADD_11602

//BasicMUL48_894 replaced by BasicMUL48_970

//BasicMUL48_895 replaced by BasicMUL48_967

//BasicMUL48_896 replaced by BasicMUL48_970

//ADD_11350 replaced by ADD_11602

//ADD_11349 replaced by ADD_11602

//ADD_11348 replaced by ADD_11602

//ADD_11353 replaced by ADD_11601

//ADD_11352 replaced by ADD_11602

//ADD_11351 replaced by ADD_11602

//ADD_11355 replaced by ADD_11602

//ADD_11354 replaced by ADD_11602

//BasicMUL48_897 replaced by BasicMUL48_971

//BasicMUL48_898 replaced by BasicMUL48_970

//BasicMUL48_899 replaced by BasicMUL48_971

//ADD_11358 replaced by ADD_11595

//ADD_11357 replaced by ADD_11602

//ADD_11356 replaced by ADD_11602

//ADD_11361 replaced by ADD_11592

//ADD_11360 replaced by ADD_11602

//ADD_11359 replaced by ADD_11602

//ADD_11364 replaced by ADD_11592

//ADD_11363 replaced by ADD_11602

//ADD_11362 replaced by ADD_11602

//ADD_11367 replaced by ADD_11595

//ADD_11366 replaced by ADD_11602

//ADD_11365 replaced by ADD_11602

//BasicMUL48_900 replaced by BasicMUL48_970

//BasicMUL48_901 replaced by BasicMUL48_967

//BasicMUL48_902 replaced by BasicMUL48_970

//ADD_11370 replaced by ADD_11563

//ADD_11369 replaced by ADD_11602

//ADD_11368 replaced by ADD_11602

//ADD_11373 replaced by ADD_11560

//ADD_11372 replaced by ADD_11602

//ADD_11371 replaced by ADD_11602

//ADD_11376 replaced by ADD_11560

//ADD_11375 replaced by ADD_11602

//ADD_11374 replaced by ADD_11602

//ADD_11379 replaced by ADD_11563

//ADD_11378 replaced by ADD_11602

//ADD_11377 replaced by ADD_11602

//BasicMUL48_903 replaced by BasicMUL48_967

//BasicMUL48_904 replaced by BasicMUL48_958

//BasicMUL48_905 replaced by BasicMUL48_967

//ADD_11382 replaced by ADD_11595

//ADD_11381 replaced by ADD_11602

//ADD_11380 replaced by ADD_11602

//ADD_11385 replaced by ADD_11592

//ADD_11384 replaced by ADD_11602

//ADD_11383 replaced by ADD_11602

//ADD_11388 replaced by ADD_11592

//ADD_11387 replaced by ADD_11602

//ADD_11386 replaced by ADD_11602

//ADD_11391 replaced by ADD_11595

//ADD_11390 replaced by ADD_11602

//ADD_11389 replaced by ADD_11602

//BasicMUL48_906 replaced by BasicMUL48_970

//BasicMUL48_907 replaced by BasicMUL48_967

//BasicMUL48_908 replaced by BasicMUL48_970

//ADD_11394 replaced by ADD_11602

//ADD_11393 replaced by ADD_11602

//ADD_11392 replaced by ADD_11602

//ADD_11397 replaced by ADD_11601

//ADD_11396 replaced by ADD_11602

//ADD_11395 replaced by ADD_11602

//ADD_11399 replaced by ADD_11602

//ADD_11398 replaced by ADD_11602

//BasicMUL48_909 replaced by BasicMUL48_971

//BasicMUL48_910 replaced by BasicMUL48_970

//BasicMUL48_911 replaced by BasicMUL48_971

//ADD_11402 replaced by ADD_11595

//ADD_11401 replaced by ADD_11602

//ADD_11400 replaced by ADD_11602

//ADD_11405 replaced by ADD_11592

//ADD_11404 replaced by ADD_11602

//ADD_11403 replaced by ADD_11602

//ADD_11408 replaced by ADD_11592

//ADD_11407 replaced by ADD_11602

//ADD_11406 replaced by ADD_11602

//ADD_11411 replaced by ADD_11595

//ADD_11410 replaced by ADD_11602

//ADD_11409 replaced by ADD_11602

//BasicMUL48_912 replaced by BasicMUL48_970

//BasicMUL48_913 replaced by BasicMUL48_967

//BasicMUL48_914 replaced by BasicMUL48_970

//ADD_11414 replaced by ADD_11602

//ADD_11413 replaced by ADD_11602

//ADD_11412 replaced by ADD_11602

//ADD_11417 replaced by ADD_11601

//ADD_11416 replaced by ADD_11602

//ADD_11415 replaced by ADD_11602

//ADD_11419 replaced by ADD_11602

//ADD_11418 replaced by ADD_11602

//BasicMUL48_915 replaced by BasicMUL48_971

//BasicMUL48_916 replaced by BasicMUL48_970

//BasicMUL48_917 replaced by BasicMUL48_971

//ADD_11422 replaced by ADD_11602

//ADD_11421 replaced by ADD_11602

//ADD_11420 replaced by ADD_11602

//ADD_11425 replaced by ADD_11601

//ADD_11424 replaced by ADD_11602

//ADD_11423 replaced by ADD_11602

//ADD_11427 replaced by ADD_11602

//ADD_11426 replaced by ADD_11602

//BasicMUL48_918 replaced by BasicMUL48_971

//BasicMUL48_919 replaced by BasicMUL48_970

//BasicMUL48_920 replaced by BasicMUL48_971

//ADD_11430 replaced by ADD_11595

//ADD_11429 replaced by ADD_11602

//ADD_11428 replaced by ADD_11602

//ADD_11433 replaced by ADD_11592

//ADD_11432 replaced by ADD_11602

//ADD_11431 replaced by ADD_11602

//ADD_11436 replaced by ADD_11592

//ADD_11435 replaced by ADD_11602

//ADD_11434 replaced by ADD_11602

//ADD_11439 replaced by ADD_11595

//ADD_11438 replaced by ADD_11602

//ADD_11437 replaced by ADD_11602

//BasicMUL48_921 replaced by BasicMUL48_970

//BasicMUL48_922 replaced by BasicMUL48_967

//BasicMUL48_923 replaced by BasicMUL48_970

//ADD_11442 replaced by ADD_11602

//ADD_11441 replaced by ADD_11602

//ADD_11440 replaced by ADD_11602

//ADD_11445 replaced by ADD_11601

//ADD_11444 replaced by ADD_11602

//ADD_11443 replaced by ADD_11602

//ADD_11447 replaced by ADD_11602

//ADD_11446 replaced by ADD_11602

//BasicMUL48_924 replaced by BasicMUL48_971

//BasicMUL48_925 replaced by BasicMUL48_970

//BasicMUL48_926 replaced by BasicMUL48_971

//ADD_11450 replaced by ADD_11595

//ADD_11449 replaced by ADD_11602

//ADD_11448 replaced by ADD_11602

//ADD_11453 replaced by ADD_11592

//ADD_11452 replaced by ADD_11602

//ADD_11451 replaced by ADD_11602

//ADD_11456 replaced by ADD_11592

//ADD_11455 replaced by ADD_11602

//ADD_11454 replaced by ADD_11602

//ADD_11459 replaced by ADD_11595

//ADD_11458 replaced by ADD_11602

//ADD_11457 replaced by ADD_11602

//BasicMUL48_927 replaced by BasicMUL48_970

//BasicMUL48_928 replaced by BasicMUL48_967

//BasicMUL48_929 replaced by BasicMUL48_970

//ADD_11462 replaced by ADD_11563

//ADD_11461 replaced by ADD_11602

//ADD_11460 replaced by ADD_11602

//ADD_11465 replaced by ADD_11560

//ADD_11464 replaced by ADD_11602

//ADD_11463 replaced by ADD_11602

//ADD_11468 replaced by ADD_11560

//ADD_11467 replaced by ADD_11602

//ADD_11466 replaced by ADD_11602

//ADD_11471 replaced by ADD_11563

//ADD_11470 replaced by ADD_11602

//ADD_11469 replaced by ADD_11602

//BasicMUL48_930 replaced by BasicMUL48_967

//BasicMUL48_931 replaced by BasicMUL48_958

//BasicMUL48_932 replaced by BasicMUL48_967

//ADD_11474 replaced by ADD_11595

//ADD_11473 replaced by ADD_11602

//ADD_11472 replaced by ADD_11602

//ADD_11477 replaced by ADD_11592

//ADD_11476 replaced by ADD_11602

//ADD_11475 replaced by ADD_11602

//ADD_11480 replaced by ADD_11592

//ADD_11479 replaced by ADD_11602

//ADD_11478 replaced by ADD_11602

//ADD_11483 replaced by ADD_11595

//ADD_11482 replaced by ADD_11602

//ADD_11481 replaced by ADD_11602

//BasicMUL48_933 replaced by BasicMUL48_970

//BasicMUL48_934 replaced by BasicMUL48_967

//BasicMUL48_935 replaced by BasicMUL48_970

//ADD_11486 replaced by ADD_11602

//ADD_11485 replaced by ADD_11602

//ADD_11484 replaced by ADD_11602

//ADD_11489 replaced by ADD_11601

//ADD_11488 replaced by ADD_11602

//ADD_11487 replaced by ADD_11602

//ADD_11491 replaced by ADD_11602

//ADD_11490 replaced by ADD_11602

//BasicMUL48_936 replaced by BasicMUL48_971

//BasicMUL48_937 replaced by BasicMUL48_970

//BasicMUL48_938 replaced by BasicMUL48_971

//ADD_11494 replaced by ADD_11595

//ADD_11493 replaced by ADD_11602

//ADD_11492 replaced by ADD_11602

//ADD_11497 replaced by ADD_11592

//ADD_11496 replaced by ADD_11602

//ADD_11495 replaced by ADD_11602

//ADD_11500 replaced by ADD_11592

//ADD_11499 replaced by ADD_11602

//ADD_11498 replaced by ADD_11602

//ADD_11503 replaced by ADD_11595

//ADD_11502 replaced by ADD_11602

//ADD_11501 replaced by ADD_11602

//BasicMUL48_939 replaced by BasicMUL48_970

//BasicMUL48_940 replaced by BasicMUL48_967

//BasicMUL48_941 replaced by BasicMUL48_970

//ADD_11506 replaced by ADD_11602

//ADD_11505 replaced by ADD_11602

//ADD_11504 replaced by ADD_11602

//ADD_11509 replaced by ADD_11601

//ADD_11508 replaced by ADD_11602

//ADD_11507 replaced by ADD_11602

//ADD_11511 replaced by ADD_11602

//ADD_11510 replaced by ADD_11602

//BasicMUL48_942 replaced by BasicMUL48_971

//BasicMUL48_943 replaced by BasicMUL48_970

//BasicMUL48_944 replaced by BasicMUL48_971

//ADD_11514 replaced by ADD_11602

//ADD_11513 replaced by ADD_11602

//ADD_11512 replaced by ADD_11602

//ADD_11517 replaced by ADD_11601

//ADD_11516 replaced by ADD_11602

//ADD_11515 replaced by ADD_11602

//ADD_11519 replaced by ADD_11602

//ADD_11518 replaced by ADD_11602

//BasicMUL48_945 replaced by BasicMUL48_971

//BasicMUL48_946 replaced by BasicMUL48_970

//BasicMUL48_947 replaced by BasicMUL48_971

//ADD_11522 replaced by ADD_11595

//ADD_11521 replaced by ADD_11602

//ADD_11520 replaced by ADD_11602

//ADD_11525 replaced by ADD_11592

//ADD_11524 replaced by ADD_11602

//ADD_11523 replaced by ADD_11602

//ADD_11528 replaced by ADD_11592

//ADD_11527 replaced by ADD_11602

//ADD_11526 replaced by ADD_11602

//ADD_11531 replaced by ADD_11595

//ADD_11530 replaced by ADD_11602

//ADD_11529 replaced by ADD_11602

//BasicMUL48_948 replaced by BasicMUL48_970

//BasicMUL48_949 replaced by BasicMUL48_967

//BasicMUL48_950 replaced by BasicMUL48_970

//ADD_11534 replaced by ADD_11602

//ADD_11533 replaced by ADD_11602

//ADD_11532 replaced by ADD_11602

//ADD_11537 replaced by ADD_11601

//ADD_11536 replaced by ADD_11602

//ADD_11535 replaced by ADD_11602

//ADD_11539 replaced by ADD_11602

//ADD_11538 replaced by ADD_11602

//BasicMUL48_951 replaced by BasicMUL48_971

//BasicMUL48_952 replaced by BasicMUL48_970

//BasicMUL48_953 replaced by BasicMUL48_971

//ADD_11542 replaced by ADD_11595

//ADD_11541 replaced by ADD_11602

//ADD_11540 replaced by ADD_11602

//ADD_11545 replaced by ADD_11592

//ADD_11544 replaced by ADD_11602

//ADD_11543 replaced by ADD_11602

//ADD_11548 replaced by ADD_11592

//ADD_11547 replaced by ADD_11602

//ADD_11546 replaced by ADD_11602

//ADD_11551 replaced by ADD_11595

//ADD_11550 replaced by ADD_11602

//ADD_11549 replaced by ADD_11602

//BasicMUL48_954 replaced by BasicMUL48_970

//BasicMUL48_955 replaced by BasicMUL48_967

//BasicMUL48_956 replaced by BasicMUL48_970

//ADD_11554 replaced by ADD_11563

//ADD_11553 replaced by ADD_11602

//ADD_11552 replaced by ADD_11602

//ADD_11557 replaced by ADD_11560

//ADD_11556 replaced by ADD_11602

//ADD_11555 replaced by ADD_11602

module ADD_11560 (
  input      [4:0]    io_A_0,
  input      [4:0]    io_A_1,
  input               io_CIN,
  output     [5:0]    io_S
);

  wire       [5:0]    _zz_io_S;
  wire       [5:0]    _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {5'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_11559 replaced by ADD_11602

//ADD_11558 replaced by ADD_11602

module ADD_11563 (
  input      [3:0]    io_A_0,
  input      [3:0]    io_A_1,
  input               io_CIN,
  output     [4:0]    io_S
);

  wire       [4:0]    _zz_io_S;
  wire       [4:0]    _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {4'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_11562 replaced by ADD_11602

//ADD_11561 replaced by ADD_11602

//BasicMUL48_957 replaced by BasicMUL48_967

module BasicMUL48_958 (
  input      [50:0]   io_a,
  input      [50:0]   io_b,
  output     [101:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [51:0]   mul_io_a;
  wire       [102:0]  mul_io_p;
  wire       [101:0]  p;

  BasicMAC48_971 mul (
    .io_a   (mul_io_a[51:0] ), //i
    .io_b   (io_b[50:0]     ), //i
    .io_c   (51'h0          ), //i
    .io_ce  (1'b1           ), //i
    .io_p   (mul_io_p[102:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  assign io_p = p;
  assign mul_io_a = {1'd0, io_a};
  assign p = mul_io_p[101:0];

endmodule

//BasicMUL48_959 replaced by BasicMUL48_967

//ADD_11566 replaced by ADD_11595

//ADD_11565 replaced by ADD_11602

//ADD_11564 replaced by ADD_11602

//ADD_11569 replaced by ADD_11592

//ADD_11568 replaced by ADD_11602

//ADD_11567 replaced by ADD_11602

//ADD_11572 replaced by ADD_11592

//ADD_11571 replaced by ADD_11602

//ADD_11570 replaced by ADD_11602

//ADD_11575 replaced by ADD_11595

//ADD_11574 replaced by ADD_11602

//ADD_11573 replaced by ADD_11602

//BasicMUL48_960 replaced by BasicMUL48_970

//BasicMUL48_961 replaced by BasicMUL48_967

//BasicMUL48_962 replaced by BasicMUL48_970

//ADD_11578 replaced by ADD_11602

//ADD_11577 replaced by ADD_11602

//ADD_11576 replaced by ADD_11602

//ADD_11581 replaced by ADD_11601

//ADD_11580 replaced by ADD_11602

//ADD_11579 replaced by ADD_11602

//ADD_11583 replaced by ADD_11602

//ADD_11582 replaced by ADD_11602

//BasicMUL48_963 replaced by BasicMUL48_971

//BasicMUL48_964 replaced by BasicMUL48_970

//BasicMUL48_965 replaced by BasicMUL48_971

//ADD_11586 replaced by ADD_11595

//ADD_11585 replaced by ADD_11602

//ADD_11584 replaced by ADD_11602

//ADD_11589 replaced by ADD_11592

//ADD_11588 replaced by ADD_11602

//ADD_11587 replaced by ADD_11602

module ADD_11592 (
  input      [2:0]    io_A_0,
  input      [2:0]    io_A_1,
  input               io_CIN,
  output     [3:0]    io_S
);

  wire       [3:0]    _zz_io_S;
  wire       [3:0]    _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {3'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_11591 replaced by ADD_11602

//ADD_11590 replaced by ADD_11602

module ADD_11595 (
  input      [1:0]    io_A_0,
  input      [1:0]    io_A_1,
  input               io_CIN,
  output     [2:0]    io_S
);

  wire       [2:0]    _zz_io_S;
  wire       [2:0]    _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {2'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_11594 replaced by ADD_11602

//ADD_11593 replaced by ADD_11602

//BasicMUL48_966 replaced by BasicMUL48_970

module BasicMUL48_967 (
  input      [49:0]   io_a,
  input      [49:0]   io_b,
  output     [99:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [51:0]   mul_io_a;
  wire       [50:0]   mul_io_b;
  wire       [102:0]  mul_io_p;
  wire       [99:0]   p;

  BasicMAC48_971 mul (
    .io_a   (mul_io_a[51:0] ), //i
    .io_b   (mul_io_b[50:0] ), //i
    .io_c   (51'h0          ), //i
    .io_ce  (1'b1           ), //i
    .io_p   (mul_io_p[102:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  assign io_p = p;
  assign mul_io_a = {2'd0, io_a};
  assign mul_io_b = {1'd0, io_b};
  assign p = mul_io_p[99:0];

endmodule

//BasicMUL48_968 replaced by BasicMUL48_970

//ADD_11598 replaced by ADD_11602

//ADD_11597 replaced by ADD_11602

//ADD_11596 replaced by ADD_11602

module ADD_11601 (
  input      [0:0]    io_A_0,
  input      [0:0]    io_A_1,
  input               io_CIN,
  output     [1:0]    io_S
);

  wire       [1:0]    _zz_io_S;
  wire       [1:0]    _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {1'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//ADD_11600 replaced by ADD_11602

//ADD_11599 replaced by ADD_11602

//ADD_11603 replaced by ADD_11602

module ADD_11602 (
  input      [47:0]   io_A_0,
  input      [47:0]   io_A_1,
  input               io_CIN,
  output     [48:0]   io_S
);

  wire       [48:0]   _zz_io_S;
  wire       [48:0]   _zz_io_S_1;
  wire       [0:0]    _zz_io_S_2;

  assign _zz_io_S = ({1'b0,io_A_0} + {1'b0,io_A_1});
  assign _zz_io_S_2 = io_CIN;
  assign _zz_io_S_1 = {48'd0, _zz_io_S_2};
  assign io_S = (_zz_io_S + _zz_io_S_1);

endmodule

//BasicMUL48_969 replaced by BasicMUL48_971

module BasicMUL48_970 (
  input      [48:0]   io_a,
  input      [48:0]   io_b,
  output     [97:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [51:0]   mul_io_a;
  wire       [50:0]   mul_io_b;
  wire       [102:0]  mul_io_p;
  wire       [97:0]   p;

  BasicMAC48_971 mul (
    .io_a   (mul_io_a[51:0] ), //i
    .io_b   (mul_io_b[50:0] ), //i
    .io_c   (51'h0          ), //i
    .io_ce  (1'b1           ), //i
    .io_p   (mul_io_p[102:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  assign io_p = p;
  assign mul_io_a = {3'd0, io_a};
  assign mul_io_b = {2'd0, io_b};
  assign p = mul_io_p[97:0];

endmodule

module BasicMUL48_971 (
  input      [47:0]   io_a,
  input      [47:0]   io_b,
  output     [95:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [51:0]   mul_io_a;
  wire       [50:0]   mul_io_b;
  wire       [102:0]  mul_io_p;
  wire       [95:0]   p;

  BasicMAC48_971 mul (
    .io_a   (mul_io_a[51:0] ), //i
    .io_b   (mul_io_b[50:0] ), //i
    .io_c   (51'h0          ), //i
    .io_ce  (1'b1           ), //i
    .io_p   (mul_io_p[102:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  assign io_p = p;
  assign mul_io_a = {4'd0, io_a};
  assign mul_io_b = {3'd0, io_b};
  assign p = mul_io_p[95:0];

endmodule

//BasicMAC48 replaced by BasicMAC48_971

//BasicMAC48_1 replaced by BasicMAC48_971

//BasicMAC48_2 replaced by BasicMAC48_971

//BasicMAC48_3 replaced by BasicMAC48_971

//BasicMAC48_4 replaced by BasicMAC48_971

//BasicMAC48_5 replaced by BasicMAC48_971

//BasicMAC48_6 replaced by BasicMAC48_971

//BasicMAC48_7 replaced by BasicMAC48_971

//BasicMAC48_8 replaced by BasicMAC48_971

//BasicMAC48_9 replaced by BasicMAC48_971

//BasicMAC48_10 replaced by BasicMAC48_971

//BasicMAC48_11 replaced by BasicMAC48_971

//BasicMAC48_12 replaced by BasicMAC48_971

//BasicMAC48_13 replaced by BasicMAC48_971

//BasicMAC48_14 replaced by BasicMAC48_971

//BasicMAC48_15 replaced by BasicMAC48_971

//BasicMAC48_16 replaced by BasicMAC48_971

//BasicMAC48_17 replaced by BasicMAC48_971

//BasicMAC48_18 replaced by BasicMAC48_971

//BasicMAC48_19 replaced by BasicMAC48_971

//BasicMAC48_20 replaced by BasicMAC48_971

//BasicMAC48_21 replaced by BasicMAC48_971

//BasicMAC48_22 replaced by BasicMAC48_971

//BasicMAC48_23 replaced by BasicMAC48_971

//BasicMAC48_24 replaced by BasicMAC48_971

//BasicMAC48_25 replaced by BasicMAC48_971

//BasicMAC48_26 replaced by BasicMAC48_971

//BasicMAC48_27 replaced by BasicMAC48_971

//BasicMAC48_28 replaced by BasicMAC48_971

//BasicMAC48_29 replaced by BasicMAC48_971

//BasicMAC48_30 replaced by BasicMAC48_971

//BasicMAC48_31 replaced by BasicMAC48_971

//BasicMAC48_32 replaced by BasicMAC48_971

//BasicMAC48_33 replaced by BasicMAC48_971

//BasicMAC48_34 replaced by BasicMAC48_971

//BasicMAC48_35 replaced by BasicMAC48_971

//BasicMAC48_36 replaced by BasicMAC48_971

//BasicMAC48_37 replaced by BasicMAC48_971

//BasicMAC48_38 replaced by BasicMAC48_971

//BasicMAC48_39 replaced by BasicMAC48_971

//BasicMAC48_40 replaced by BasicMAC48_971

//BasicMAC48_41 replaced by BasicMAC48_971

//BasicMAC48_42 replaced by BasicMAC48_971

//BasicMAC48_43 replaced by BasicMAC48_971

//BasicMAC48_44 replaced by BasicMAC48_971

//BasicMAC48_45 replaced by BasicMAC48_971

//BasicMAC48_46 replaced by BasicMAC48_971

//BasicMAC48_47 replaced by BasicMAC48_971

//BasicMAC48_48 replaced by BasicMAC48_971

//BasicMAC48_49 replaced by BasicMAC48_971

//BasicMAC48_50 replaced by BasicMAC48_971

//BasicMAC48_51 replaced by BasicMAC48_971

//BasicMAC48_52 replaced by BasicMAC48_971

//BasicMAC48_53 replaced by BasicMAC48_971

//BasicMAC48_54 replaced by BasicMAC48_971

//BasicMAC48_55 replaced by BasicMAC48_971

//BasicMAC48_56 replaced by BasicMAC48_971

//BasicMAC48_57 replaced by BasicMAC48_971

//BasicMAC48_58 replaced by BasicMAC48_971

//BasicMAC48_59 replaced by BasicMAC48_971

//BasicMAC48_60 replaced by BasicMAC48_971

//BasicMAC48_61 replaced by BasicMAC48_971

//BasicMAC48_62 replaced by BasicMAC48_971

//BasicMAC48_63 replaced by BasicMAC48_971

//BasicMAC48_64 replaced by BasicMAC48_971

//BasicMAC48_65 replaced by BasicMAC48_971

//BasicMAC48_66 replaced by BasicMAC48_971

//BasicMAC48_67 replaced by BasicMAC48_971

//BasicMAC48_68 replaced by BasicMAC48_971

//BasicMAC48_69 replaced by BasicMAC48_971

//BasicMAC48_70 replaced by BasicMAC48_971

//BasicMAC48_71 replaced by BasicMAC48_971

//BasicMAC48_72 replaced by BasicMAC48_971

//BasicMAC48_73 replaced by BasicMAC48_971

//BasicMAC48_74 replaced by BasicMAC48_971

//BasicMAC48_75 replaced by BasicMAC48_971

//BasicMAC48_76 replaced by BasicMAC48_971

//BasicMAC48_77 replaced by BasicMAC48_971

//BasicMAC48_78 replaced by BasicMAC48_971

//BasicMAC48_79 replaced by BasicMAC48_971

//BasicMAC48_80 replaced by BasicMAC48_971

//BasicMAC48_81 replaced by BasicMAC48_971

//BasicMAC48_82 replaced by BasicMAC48_971

//BasicMAC48_83 replaced by BasicMAC48_971

//BasicMAC48_84 replaced by BasicMAC48_971

//BasicMAC48_85 replaced by BasicMAC48_971

//BasicMAC48_86 replaced by BasicMAC48_971

//BasicMAC48_87 replaced by BasicMAC48_971

//BasicMAC48_88 replaced by BasicMAC48_971

//BasicMAC48_89 replaced by BasicMAC48_971

//BasicMAC48_90 replaced by BasicMAC48_971

//BasicMAC48_91 replaced by BasicMAC48_971

//BasicMAC48_92 replaced by BasicMAC48_971

//BasicMAC48_93 replaced by BasicMAC48_971

//BasicMAC48_94 replaced by BasicMAC48_971

//BasicMAC48_95 replaced by BasicMAC48_971

//BasicMAC48_96 replaced by BasicMAC48_971

//BasicMAC48_97 replaced by BasicMAC48_971

//BasicMAC48_98 replaced by BasicMAC48_971

//BasicMAC48_99 replaced by BasicMAC48_971

//BasicMAC48_100 replaced by BasicMAC48_971

//BasicMAC48_101 replaced by BasicMAC48_971

//BasicMAC48_102 replaced by BasicMAC48_971

//BasicMAC48_103 replaced by BasicMAC48_971

//BasicMAC48_104 replaced by BasicMAC48_971

//BasicMAC48_105 replaced by BasicMAC48_971

//BasicMAC48_106 replaced by BasicMAC48_971

//BasicMAC48_107 replaced by BasicMAC48_971

//BasicMAC48_108 replaced by BasicMAC48_971

//BasicMAC48_109 replaced by BasicMAC48_971

//BasicMAC48_110 replaced by BasicMAC48_971

//BasicMAC48_111 replaced by BasicMAC48_971

//BasicMAC48_112 replaced by BasicMAC48_971

//BasicMAC48_113 replaced by BasicMAC48_971

//BasicMAC48_114 replaced by BasicMAC48_971

//BasicMAC48_115 replaced by BasicMAC48_971

//BasicMAC48_116 replaced by BasicMAC48_971

//BasicMAC48_117 replaced by BasicMAC48_971

//BasicMAC48_118 replaced by BasicMAC48_971

//BasicMAC48_119 replaced by BasicMAC48_971

//BasicMAC48_120 replaced by BasicMAC48_971

//BasicMAC48_121 replaced by BasicMAC48_971

//BasicMAC48_122 replaced by BasicMAC48_971

//BasicMAC48_123 replaced by BasicMAC48_971

//BasicMAC48_124 replaced by BasicMAC48_971

//BasicMAC48_125 replaced by BasicMAC48_971

//BasicMAC48_126 replaced by BasicMAC48_971

//BasicMAC48_127 replaced by BasicMAC48_971

//BasicMAC48_128 replaced by BasicMAC48_971

//BasicMAC48_129 replaced by BasicMAC48_971

//BasicMAC48_130 replaced by BasicMAC48_971

//BasicMAC48_131 replaced by BasicMAC48_971

//BasicMAC48_132 replaced by BasicMAC48_971

//BasicMAC48_133 replaced by BasicMAC48_971

//BasicMAC48_134 replaced by BasicMAC48_971

//BasicMAC48_135 replaced by BasicMAC48_971

//BasicMAC48_136 replaced by BasicMAC48_971

//BasicMAC48_137 replaced by BasicMAC48_971

//BasicMAC48_138 replaced by BasicMAC48_971

//BasicMAC48_139 replaced by BasicMAC48_971

//BasicMAC48_140 replaced by BasicMAC48_971

//BasicMAC48_141 replaced by BasicMAC48_971

//BasicMAC48_142 replaced by BasicMAC48_971

//BasicMAC48_143 replaced by BasicMAC48_971

//BasicMAC48_144 replaced by BasicMAC48_971

//BasicMAC48_145 replaced by BasicMAC48_971

//BasicMAC48_146 replaced by BasicMAC48_971

//BasicMAC48_147 replaced by BasicMAC48_971

//BasicMAC48_148 replaced by BasicMAC48_971

//BasicMAC48_149 replaced by BasicMAC48_971

//BasicMAC48_150 replaced by BasicMAC48_971

//BasicMAC48_151 replaced by BasicMAC48_971

//BasicMAC48_152 replaced by BasicMAC48_971

//BasicMAC48_153 replaced by BasicMAC48_971

//BasicMAC48_154 replaced by BasicMAC48_971

//BasicMAC48_155 replaced by BasicMAC48_971

//BasicMAC48_156 replaced by BasicMAC48_971

//BasicMAC48_157 replaced by BasicMAC48_971

//BasicMAC48_158 replaced by BasicMAC48_971

//BasicMAC48_159 replaced by BasicMAC48_971

//BasicMAC48_160 replaced by BasicMAC48_971

//BasicMAC48_161 replaced by BasicMAC48_971

//BasicMAC48_162 replaced by BasicMAC48_971

//BasicMAC48_163 replaced by BasicMAC48_971

//BasicMAC48_164 replaced by BasicMAC48_971

//BasicMAC48_165 replaced by BasicMAC48_971

//BasicMAC48_166 replaced by BasicMAC48_971

//BasicMAC48_167 replaced by BasicMAC48_971

//BasicMAC48_168 replaced by BasicMAC48_971

//BasicMAC48_169 replaced by BasicMAC48_971

//BasicMAC48_170 replaced by BasicMAC48_971

//BasicMAC48_171 replaced by BasicMAC48_971

//BasicMAC48_172 replaced by BasicMAC48_971

//BasicMAC48_173 replaced by BasicMAC48_971

//BasicMAC48_174 replaced by BasicMAC48_971

//BasicMAC48_175 replaced by BasicMAC48_971

//BasicMAC48_176 replaced by BasicMAC48_971

//BasicMAC48_177 replaced by BasicMAC48_971

//BasicMAC48_178 replaced by BasicMAC48_971

//BasicMAC48_179 replaced by BasicMAC48_971

//BasicMAC48_180 replaced by BasicMAC48_971

//BasicMAC48_181 replaced by BasicMAC48_971

//BasicMAC48_182 replaced by BasicMAC48_971

//BasicMAC48_183 replaced by BasicMAC48_971

//BasicMAC48_184 replaced by BasicMAC48_971

//BasicMAC48_185 replaced by BasicMAC48_971

//BasicMAC48_186 replaced by BasicMAC48_971

//BasicMAC48_187 replaced by BasicMAC48_971

//BasicMAC48_188 replaced by BasicMAC48_971

//BasicMAC48_189 replaced by BasicMAC48_971

//BasicMAC48_190 replaced by BasicMAC48_971

//BasicMAC48_191 replaced by BasicMAC48_971

//BasicMAC48_192 replaced by BasicMAC48_971

//BasicMAC48_193 replaced by BasicMAC48_971

//BasicMAC48_194 replaced by BasicMAC48_971

//BasicMAC48_195 replaced by BasicMAC48_971

//BasicMAC48_196 replaced by BasicMAC48_971

//BasicMAC48_197 replaced by BasicMAC48_971

//BasicMAC48_198 replaced by BasicMAC48_971

//BasicMAC48_199 replaced by BasicMAC48_971

//BasicMAC48_200 replaced by BasicMAC48_971

//BasicMAC48_201 replaced by BasicMAC48_971

//BasicMAC48_202 replaced by BasicMAC48_971

//BasicMAC48_203 replaced by BasicMAC48_971

//BasicMAC48_204 replaced by BasicMAC48_971

//BasicMAC48_205 replaced by BasicMAC48_971

//BasicMAC48_206 replaced by BasicMAC48_971

//BasicMAC48_207 replaced by BasicMAC48_971

//BasicMAC48_208 replaced by BasicMAC48_971

//BasicMAC48_209 replaced by BasicMAC48_971

//BasicMAC48_210 replaced by BasicMAC48_971

//BasicMAC48_211 replaced by BasicMAC48_971

//BasicMAC48_212 replaced by BasicMAC48_971

//BasicMAC48_213 replaced by BasicMAC48_971

//BasicMAC48_214 replaced by BasicMAC48_971

//BasicMAC48_215 replaced by BasicMAC48_971

//BasicMAC48_216 replaced by BasicMAC48_971

//BasicMAC48_217 replaced by BasicMAC48_971

//BasicMAC48_218 replaced by BasicMAC48_971

//BasicMAC48_219 replaced by BasicMAC48_971

//BasicMAC48_220 replaced by BasicMAC48_971

//BasicMAC48_221 replaced by BasicMAC48_971

//BasicMAC48_222 replaced by BasicMAC48_971

//BasicMAC48_223 replaced by BasicMAC48_971

//BasicMAC48_224 replaced by BasicMAC48_971

//BasicMAC48_225 replaced by BasicMAC48_971

//BasicMAC48_226 replaced by BasicMAC48_971

//BasicMAC48_227 replaced by BasicMAC48_971

//BasicMAC48_228 replaced by BasicMAC48_971

//BasicMAC48_229 replaced by BasicMAC48_971

//BasicMAC48_230 replaced by BasicMAC48_971

//BasicMAC48_231 replaced by BasicMAC48_971

//BasicMAC48_232 replaced by BasicMAC48_971

//BasicMAC48_233 replaced by BasicMAC48_971

//BasicMAC48_234 replaced by BasicMAC48_971

//BasicMAC48_235 replaced by BasicMAC48_971

//BasicMAC48_236 replaced by BasicMAC48_971

//BasicMAC48_237 replaced by BasicMAC48_971

//BasicMAC48_238 replaced by BasicMAC48_971

//BasicMAC48_239 replaced by BasicMAC48_971

//BasicMAC48_240 replaced by BasicMAC48_971

//BasicMAC48_241 replaced by BasicMAC48_971

//BasicMAC48_242 replaced by BasicMAC48_971

//BasicMAC48_243 replaced by BasicMAC48_971

//BasicMAC48_244 replaced by BasicMAC48_971

//BasicMAC48_245 replaced by BasicMAC48_971

//BasicMAC48_246 replaced by BasicMAC48_971

//BasicMAC48_247 replaced by BasicMAC48_971

//BasicMAC48_248 replaced by BasicMAC48_971

//BasicMAC48_249 replaced by BasicMAC48_971

//BasicMAC48_250 replaced by BasicMAC48_971

//BasicMAC48_251 replaced by BasicMAC48_971

//BasicMAC48_252 replaced by BasicMAC48_971

//BasicMAC48_253 replaced by BasicMAC48_971

//BasicMAC48_254 replaced by BasicMAC48_971

//BasicMAC48_255 replaced by BasicMAC48_971

//BasicMAC48_256 replaced by BasicMAC48_971

//BasicMAC48_257 replaced by BasicMAC48_971

//BasicMAC48_258 replaced by BasicMAC48_971

//BasicMAC48_259 replaced by BasicMAC48_971

//BasicMAC48_260 replaced by BasicMAC48_971

//BasicMAC48_261 replaced by BasicMAC48_971

//BasicMAC48_262 replaced by BasicMAC48_971

//BasicMAC48_263 replaced by BasicMAC48_971

//BasicMAC48_264 replaced by BasicMAC48_971

//BasicMAC48_265 replaced by BasicMAC48_971

//BasicMAC48_266 replaced by BasicMAC48_971

//BasicMAC48_267 replaced by BasicMAC48_971

//BasicMAC48_268 replaced by BasicMAC48_971

//BasicMAC48_269 replaced by BasicMAC48_971

//BasicMAC48_270 replaced by BasicMAC48_971

//BasicMAC48_271 replaced by BasicMAC48_971

//BasicMAC48_272 replaced by BasicMAC48_971

//BasicMAC48_273 replaced by BasicMAC48_971

//BasicMAC48_274 replaced by BasicMAC48_971

//BasicMAC48_275 replaced by BasicMAC48_971

//BasicMAC48_276 replaced by BasicMAC48_971

//BasicMAC48_277 replaced by BasicMAC48_971

//BasicMAC48_278 replaced by BasicMAC48_971

//BasicMAC48_279 replaced by BasicMAC48_971

//BasicMAC48_280 replaced by BasicMAC48_971

//BasicMAC48_281 replaced by BasicMAC48_971

//BasicMAC48_282 replaced by BasicMAC48_971

//BasicMAC48_283 replaced by BasicMAC48_971

//BasicMAC48_284 replaced by BasicMAC48_971

//BasicMAC48_285 replaced by BasicMAC48_971

//BasicMAC48_286 replaced by BasicMAC48_971

//BasicMAC48_287 replaced by BasicMAC48_971

//BasicMAC48_288 replaced by BasicMAC48_971

//BasicMAC48_289 replaced by BasicMAC48_971

//BasicMAC48_290 replaced by BasicMAC48_971

//BasicMAC48_291 replaced by BasicMAC48_971

//BasicMAC48_292 replaced by BasicMAC48_971

//BasicMAC48_293 replaced by BasicMAC48_971

//BasicMAC48_294 replaced by BasicMAC48_971

//BasicMAC48_295 replaced by BasicMAC48_971

//BasicMAC48_296 replaced by BasicMAC48_971

//BasicMAC48_297 replaced by BasicMAC48_971

//BasicMAC48_298 replaced by BasicMAC48_971

//BasicMAC48_299 replaced by BasicMAC48_971

//BasicMAC48_300 replaced by BasicMAC48_971

//BasicMAC48_301 replaced by BasicMAC48_971

//BasicMAC48_302 replaced by BasicMAC48_971

//BasicMAC48_303 replaced by BasicMAC48_971

//BasicMAC48_304 replaced by BasicMAC48_971

//BasicMAC48_305 replaced by BasicMAC48_971

//BasicMAC48_306 replaced by BasicMAC48_971

//BasicMAC48_307 replaced by BasicMAC48_971

//BasicMAC48_308 replaced by BasicMAC48_971

//BasicMAC48_309 replaced by BasicMAC48_971

//BasicMAC48_310 replaced by BasicMAC48_971

//BasicMAC48_311 replaced by BasicMAC48_971

//BasicMAC48_312 replaced by BasicMAC48_971

//BasicMAC48_313 replaced by BasicMAC48_971

//BasicMAC48_314 replaced by BasicMAC48_971

//BasicMAC48_315 replaced by BasicMAC48_971

//BasicMAC48_316 replaced by BasicMAC48_971

//BasicMAC48_317 replaced by BasicMAC48_971

//BasicMAC48_318 replaced by BasicMAC48_971

//BasicMAC48_319 replaced by BasicMAC48_971

//BasicMAC48_320 replaced by BasicMAC48_971

//BasicMAC48_321 replaced by BasicMAC48_971

//BasicMAC48_322 replaced by BasicMAC48_971

//BasicMAC48_323 replaced by BasicMAC48_971

//BasicMAC48_324 replaced by BasicMAC48_971

//BasicMAC48_325 replaced by BasicMAC48_971

//BasicMAC48_326 replaced by BasicMAC48_971

//BasicMAC48_327 replaced by BasicMAC48_971

//BasicMAC48_328 replaced by BasicMAC48_971

//BasicMAC48_329 replaced by BasicMAC48_971

//BasicMAC48_330 replaced by BasicMAC48_971

//BasicMAC48_331 replaced by BasicMAC48_971

//BasicMAC48_332 replaced by BasicMAC48_971

//BasicMAC48_333 replaced by BasicMAC48_971

//BasicMAC48_334 replaced by BasicMAC48_971

//BasicMAC48_335 replaced by BasicMAC48_971

//BasicMAC48_336 replaced by BasicMAC48_971

//BasicMAC48_337 replaced by BasicMAC48_971

//BasicMAC48_338 replaced by BasicMAC48_971

//BasicMAC48_339 replaced by BasicMAC48_971

//BasicMAC48_340 replaced by BasicMAC48_971

//BasicMAC48_341 replaced by BasicMAC48_971

//BasicMAC48_342 replaced by BasicMAC48_971

//BasicMAC48_343 replaced by BasicMAC48_971

//BasicMAC48_344 replaced by BasicMAC48_971

//BasicMAC48_345 replaced by BasicMAC48_971

//BasicMAC48_346 replaced by BasicMAC48_971

//BasicMAC48_347 replaced by BasicMAC48_971

//BasicMAC48_348 replaced by BasicMAC48_971

//BasicMAC48_349 replaced by BasicMAC48_971

//BasicMAC48_350 replaced by BasicMAC48_971

//BasicMAC48_351 replaced by BasicMAC48_971

//BasicMAC48_352 replaced by BasicMAC48_971

//BasicMAC48_353 replaced by BasicMAC48_971

//BasicMAC48_354 replaced by BasicMAC48_971

//BasicMAC48_355 replaced by BasicMAC48_971

//BasicMAC48_356 replaced by BasicMAC48_971

//BasicMAC48_357 replaced by BasicMAC48_971

//BasicMAC48_358 replaced by BasicMAC48_971

//BasicMAC48_359 replaced by BasicMAC48_971

//BasicMAC48_360 replaced by BasicMAC48_971

//BasicMAC48_361 replaced by BasicMAC48_971

//BasicMAC48_362 replaced by BasicMAC48_971

//BasicMAC48_363 replaced by BasicMAC48_971

//BasicMAC48_364 replaced by BasicMAC48_971

//BasicMAC48_365 replaced by BasicMAC48_971

//BasicMAC48_366 replaced by BasicMAC48_971

//BasicMAC48_367 replaced by BasicMAC48_971

//BasicMAC48_368 replaced by BasicMAC48_971

//BasicMAC48_369 replaced by BasicMAC48_971

//BasicMAC48_370 replaced by BasicMAC48_971

//BasicMAC48_371 replaced by BasicMAC48_971

//BasicMAC48_372 replaced by BasicMAC48_971

//BasicMAC48_373 replaced by BasicMAC48_971

//BasicMAC48_374 replaced by BasicMAC48_971

//BasicMAC48_375 replaced by BasicMAC48_971

//BasicMAC48_376 replaced by BasicMAC48_971

//BasicMAC48_377 replaced by BasicMAC48_971

//BasicMAC48_378 replaced by BasicMAC48_971

//BasicMAC48_379 replaced by BasicMAC48_971

//BasicMAC48_380 replaced by BasicMAC48_971

//BasicMAC48_381 replaced by BasicMAC48_971

//BasicMAC48_382 replaced by BasicMAC48_971

//BasicMAC48_383 replaced by BasicMAC48_971

//BasicMAC48_384 replaced by BasicMAC48_971

//BasicMAC48_385 replaced by BasicMAC48_971

//BasicMAC48_386 replaced by BasicMAC48_971

//BasicMAC48_387 replaced by BasicMAC48_971

//BasicMAC48_388 replaced by BasicMAC48_971

//BasicMAC48_389 replaced by BasicMAC48_971

//BasicMAC48_390 replaced by BasicMAC48_971

//BasicMAC48_391 replaced by BasicMAC48_971

//BasicMAC48_392 replaced by BasicMAC48_971

//BasicMAC48_393 replaced by BasicMAC48_971

//BasicMAC48_394 replaced by BasicMAC48_971

//BasicMAC48_395 replaced by BasicMAC48_971

//BasicMAC48_396 replaced by BasicMAC48_971

//BasicMAC48_397 replaced by BasicMAC48_971

//BasicMAC48_398 replaced by BasicMAC48_971

//BasicMAC48_399 replaced by BasicMAC48_971

//BasicMAC48_400 replaced by BasicMAC48_971

//BasicMAC48_401 replaced by BasicMAC48_971

//BasicMAC48_402 replaced by BasicMAC48_971

//BasicMAC48_403 replaced by BasicMAC48_971

//BasicMAC48_404 replaced by BasicMAC48_971

//BasicMAC48_405 replaced by BasicMAC48_971

//BasicMAC48_406 replaced by BasicMAC48_971

//BasicMAC48_407 replaced by BasicMAC48_971

//BasicMAC48_408 replaced by BasicMAC48_971

//BasicMAC48_409 replaced by BasicMAC48_971

//BasicMAC48_410 replaced by BasicMAC48_971

//BasicMAC48_411 replaced by BasicMAC48_971

//BasicMAC48_412 replaced by BasicMAC48_971

//BasicMAC48_413 replaced by BasicMAC48_971

//BasicMAC48_414 replaced by BasicMAC48_971

//BasicMAC48_415 replaced by BasicMAC48_971

//BasicMAC48_416 replaced by BasicMAC48_971

//BasicMAC48_417 replaced by BasicMAC48_971

//BasicMAC48_418 replaced by BasicMAC48_971

//BasicMAC48_419 replaced by BasicMAC48_971

//BasicMAC48_420 replaced by BasicMAC48_971

//BasicMAC48_421 replaced by BasicMAC48_971

//BasicMAC48_422 replaced by BasicMAC48_971

//BasicMAC48_423 replaced by BasicMAC48_971

//BasicMAC48_424 replaced by BasicMAC48_971

//BasicMAC48_425 replaced by BasicMAC48_971

//BasicMAC48_426 replaced by BasicMAC48_971

//BasicMAC48_427 replaced by BasicMAC48_971

//BasicMAC48_428 replaced by BasicMAC48_971

//BasicMAC48_429 replaced by BasicMAC48_971

//BasicMAC48_430 replaced by BasicMAC48_971

//BasicMAC48_431 replaced by BasicMAC48_971

//BasicMAC48_432 replaced by BasicMAC48_971

//BasicMAC48_433 replaced by BasicMAC48_971

//BasicMAC48_434 replaced by BasicMAC48_971

//BasicMAC48_435 replaced by BasicMAC48_971

//BasicMAC48_436 replaced by BasicMAC48_971

//BasicMAC48_437 replaced by BasicMAC48_971

//BasicMAC48_438 replaced by BasicMAC48_971

//BasicMAC48_439 replaced by BasicMAC48_971

//BasicMAC48_440 replaced by BasicMAC48_971

//BasicMAC48_441 replaced by BasicMAC48_971

//BasicMAC48_442 replaced by BasicMAC48_971

//BasicMAC48_443 replaced by BasicMAC48_971

//BasicMAC48_444 replaced by BasicMAC48_971

//BasicMAC48_445 replaced by BasicMAC48_971

//BasicMAC48_446 replaced by BasicMAC48_971

//BasicMAC48_447 replaced by BasicMAC48_971

//BasicMAC48_448 replaced by BasicMAC48_971

//BasicMAC48_449 replaced by BasicMAC48_971

//BasicMAC48_450 replaced by BasicMAC48_971

//BasicMAC48_451 replaced by BasicMAC48_971

//BasicMAC48_452 replaced by BasicMAC48_971

//BasicMAC48_453 replaced by BasicMAC48_971

//BasicMAC48_454 replaced by BasicMAC48_971

//BasicMAC48_455 replaced by BasicMAC48_971

//BasicMAC48_456 replaced by BasicMAC48_971

//BasicMAC48_457 replaced by BasicMAC48_971

//BasicMAC48_458 replaced by BasicMAC48_971

//BasicMAC48_459 replaced by BasicMAC48_971

//BasicMAC48_460 replaced by BasicMAC48_971

//BasicMAC48_461 replaced by BasicMAC48_971

//BasicMAC48_462 replaced by BasicMAC48_971

//BasicMAC48_463 replaced by BasicMAC48_971

//BasicMAC48_464 replaced by BasicMAC48_971

//BasicMAC48_465 replaced by BasicMAC48_971

//BasicMAC48_466 replaced by BasicMAC48_971

//BasicMAC48_467 replaced by BasicMAC48_971

//BasicMAC48_468 replaced by BasicMAC48_971

//BasicMAC48_469 replaced by BasicMAC48_971

//BasicMAC48_470 replaced by BasicMAC48_971

//BasicMAC48_471 replaced by BasicMAC48_971

//BasicMAC48_472 replaced by BasicMAC48_971

//BasicMAC48_473 replaced by BasicMAC48_971

//BasicMAC48_474 replaced by BasicMAC48_971

//BasicMAC48_475 replaced by BasicMAC48_971

//BasicMAC48_476 replaced by BasicMAC48_971

//BasicMAC48_477 replaced by BasicMAC48_971

//BasicMAC48_478 replaced by BasicMAC48_971

//BasicMAC48_479 replaced by BasicMAC48_971

//BasicMAC48_480 replaced by BasicMAC48_971

//BasicMAC48_481 replaced by BasicMAC48_971

//BasicMAC48_482 replaced by BasicMAC48_971

//BasicMAC48_483 replaced by BasicMAC48_971

//BasicMAC48_484 replaced by BasicMAC48_971

//BasicMAC48_485 replaced by BasicMAC48_971

//BasicMAC48_486 replaced by BasicMAC48_971

//BasicMAC48_487 replaced by BasicMAC48_971

//BasicMAC48_488 replaced by BasicMAC48_971

//BasicMAC48_489 replaced by BasicMAC48_971

//BasicMAC48_490 replaced by BasicMAC48_971

//BasicMAC48_491 replaced by BasicMAC48_971

//BasicMAC48_492 replaced by BasicMAC48_971

//BasicMAC48_493 replaced by BasicMAC48_971

//BasicMAC48_494 replaced by BasicMAC48_971

//BasicMAC48_495 replaced by BasicMAC48_971

//BasicMAC48_496 replaced by BasicMAC48_971

//BasicMAC48_497 replaced by BasicMAC48_971

//BasicMAC48_498 replaced by BasicMAC48_971

//BasicMAC48_499 replaced by BasicMAC48_971

//BasicMAC48_500 replaced by BasicMAC48_971

//BasicMAC48_501 replaced by BasicMAC48_971

//BasicMAC48_502 replaced by BasicMAC48_971

//BasicMAC48_503 replaced by BasicMAC48_971

//BasicMAC48_504 replaced by BasicMAC48_971

//BasicMAC48_505 replaced by BasicMAC48_971

//BasicMAC48_506 replaced by BasicMAC48_971

//BasicMAC48_507 replaced by BasicMAC48_971

//BasicMAC48_508 replaced by BasicMAC48_971

//BasicMAC48_509 replaced by BasicMAC48_971

//BasicMAC48_510 replaced by BasicMAC48_971

//BasicMAC48_511 replaced by BasicMAC48_971

//BasicMAC48_512 replaced by BasicMAC48_971

//BasicMAC48_513 replaced by BasicMAC48_971

//BasicMAC48_514 replaced by BasicMAC48_971

//BasicMAC48_515 replaced by BasicMAC48_971

//BasicMAC48_516 replaced by BasicMAC48_971

//BasicMAC48_517 replaced by BasicMAC48_971

//BasicMAC48_518 replaced by BasicMAC48_971

//BasicMAC48_519 replaced by BasicMAC48_971

//BasicMAC48_520 replaced by BasicMAC48_971

//BasicMAC48_521 replaced by BasicMAC48_971

//BasicMAC48_522 replaced by BasicMAC48_971

//BasicMAC48_523 replaced by BasicMAC48_971

//BasicMAC48_524 replaced by BasicMAC48_971

//BasicMAC48_525 replaced by BasicMAC48_971

//BasicMAC48_526 replaced by BasicMAC48_971

//BasicMAC48_527 replaced by BasicMAC48_971

//BasicMAC48_528 replaced by BasicMAC48_971

//BasicMAC48_529 replaced by BasicMAC48_971

//BasicMAC48_530 replaced by BasicMAC48_971

//BasicMAC48_531 replaced by BasicMAC48_971

//BasicMAC48_532 replaced by BasicMAC48_971

//BasicMAC48_533 replaced by BasicMAC48_971

//BasicMAC48_534 replaced by BasicMAC48_971

//BasicMAC48_535 replaced by BasicMAC48_971

//BasicMAC48_536 replaced by BasicMAC48_971

//BasicMAC48_537 replaced by BasicMAC48_971

//BasicMAC48_538 replaced by BasicMAC48_971

//BasicMAC48_539 replaced by BasicMAC48_971

//BasicMAC48_540 replaced by BasicMAC48_971

//BasicMAC48_541 replaced by BasicMAC48_971

//BasicMAC48_542 replaced by BasicMAC48_971

//BasicMAC48_543 replaced by BasicMAC48_971

//BasicMAC48_544 replaced by BasicMAC48_971

//BasicMAC48_545 replaced by BasicMAC48_971

//BasicMAC48_546 replaced by BasicMAC48_971

//BasicMAC48_547 replaced by BasicMAC48_971

//BasicMAC48_548 replaced by BasicMAC48_971

//BasicMAC48_549 replaced by BasicMAC48_971

//BasicMAC48_550 replaced by BasicMAC48_971

//BasicMAC48_551 replaced by BasicMAC48_971

//BasicMAC48_552 replaced by BasicMAC48_971

//BasicMAC48_553 replaced by BasicMAC48_971

//BasicMAC48_554 replaced by BasicMAC48_971

//BasicMAC48_555 replaced by BasicMAC48_971

//BasicMAC48_556 replaced by BasicMAC48_971

//BasicMAC48_557 replaced by BasicMAC48_971

//BasicMAC48_558 replaced by BasicMAC48_971

//BasicMAC48_559 replaced by BasicMAC48_971

//BasicMAC48_560 replaced by BasicMAC48_971

//BasicMAC48_561 replaced by BasicMAC48_971

//BasicMAC48_562 replaced by BasicMAC48_971

//BasicMAC48_563 replaced by BasicMAC48_971

//BasicMAC48_564 replaced by BasicMAC48_971

//BasicMAC48_565 replaced by BasicMAC48_971

//BasicMAC48_566 replaced by BasicMAC48_971

//BasicMAC48_567 replaced by BasicMAC48_971

//BasicMAC48_568 replaced by BasicMAC48_971

//BasicMAC48_569 replaced by BasicMAC48_971

//BasicMAC48_570 replaced by BasicMAC48_971

//BasicMAC48_571 replaced by BasicMAC48_971

//BasicMAC48_572 replaced by BasicMAC48_971

//BasicMAC48_573 replaced by BasicMAC48_971

//BasicMAC48_574 replaced by BasicMAC48_971

//BasicMAC48_575 replaced by BasicMAC48_971

//BasicMAC48_576 replaced by BasicMAC48_971

//BasicMAC48_577 replaced by BasicMAC48_971

//BasicMAC48_578 replaced by BasicMAC48_971

//BasicMAC48_579 replaced by BasicMAC48_971

//BasicMAC48_580 replaced by BasicMAC48_971

//BasicMAC48_581 replaced by BasicMAC48_971

//BasicMAC48_582 replaced by BasicMAC48_971

//BasicMAC48_583 replaced by BasicMAC48_971

//BasicMAC48_584 replaced by BasicMAC48_971

//BasicMAC48_585 replaced by BasicMAC48_971

//BasicMAC48_586 replaced by BasicMAC48_971

//BasicMAC48_587 replaced by BasicMAC48_971

//BasicMAC48_588 replaced by BasicMAC48_971

//BasicMAC48_589 replaced by BasicMAC48_971

//BasicMAC48_590 replaced by BasicMAC48_971

//BasicMAC48_591 replaced by BasicMAC48_971

//BasicMAC48_592 replaced by BasicMAC48_971

//BasicMAC48_593 replaced by BasicMAC48_971

//BasicMAC48_594 replaced by BasicMAC48_971

//BasicMAC48_595 replaced by BasicMAC48_971

//BasicMAC48_596 replaced by BasicMAC48_971

//BasicMAC48_597 replaced by BasicMAC48_971

//BasicMAC48_598 replaced by BasicMAC48_971

//BasicMAC48_599 replaced by BasicMAC48_971

//BasicMAC48_600 replaced by BasicMAC48_971

//BasicMAC48_601 replaced by BasicMAC48_971

//BasicMAC48_602 replaced by BasicMAC48_971

//BasicMAC48_603 replaced by BasicMAC48_971

//BasicMAC48_604 replaced by BasicMAC48_971

//BasicMAC48_605 replaced by BasicMAC48_971

//BasicMAC48_606 replaced by BasicMAC48_971

//BasicMAC48_607 replaced by BasicMAC48_971

//BasicMAC48_608 replaced by BasicMAC48_971

//BasicMAC48_609 replaced by BasicMAC48_971

//BasicMAC48_610 replaced by BasicMAC48_971

//BasicMAC48_611 replaced by BasicMAC48_971

//BasicMAC48_612 replaced by BasicMAC48_971

//BasicMAC48_613 replaced by BasicMAC48_971

//BasicMAC48_614 replaced by BasicMAC48_971

//BasicMAC48_615 replaced by BasicMAC48_971

//BasicMAC48_616 replaced by BasicMAC48_971

//BasicMAC48_617 replaced by BasicMAC48_971

//BasicMAC48_618 replaced by BasicMAC48_971

//BasicMAC48_619 replaced by BasicMAC48_971

//BasicMAC48_620 replaced by BasicMAC48_971

//BasicMAC48_621 replaced by BasicMAC48_971

//BasicMAC48_622 replaced by BasicMAC48_971

//BasicMAC48_623 replaced by BasicMAC48_971

//BasicMAC48_624 replaced by BasicMAC48_971

//BasicMAC48_625 replaced by BasicMAC48_971

//BasicMAC48_626 replaced by BasicMAC48_971

//BasicMAC48_627 replaced by BasicMAC48_971

//BasicMAC48_628 replaced by BasicMAC48_971

//BasicMAC48_629 replaced by BasicMAC48_971

//BasicMAC48_630 replaced by BasicMAC48_971

//BasicMAC48_631 replaced by BasicMAC48_971

//BasicMAC48_632 replaced by BasicMAC48_971

//BasicMAC48_633 replaced by BasicMAC48_971

//BasicMAC48_634 replaced by BasicMAC48_971

//BasicMAC48_635 replaced by BasicMAC48_971

//BasicMAC48_636 replaced by BasicMAC48_971

//BasicMAC48_637 replaced by BasicMAC48_971

//BasicMAC48_638 replaced by BasicMAC48_971

//BasicMAC48_639 replaced by BasicMAC48_971

//BasicMAC48_640 replaced by BasicMAC48_971

//BasicMAC48_641 replaced by BasicMAC48_971

//BasicMAC48_642 replaced by BasicMAC48_971

//BasicMAC48_643 replaced by BasicMAC48_971

//BasicMAC48_644 replaced by BasicMAC48_971

//BasicMAC48_645 replaced by BasicMAC48_971

//BasicMAC48_646 replaced by BasicMAC48_971

//BasicMAC48_647 replaced by BasicMAC48_971

//BasicMAC48_648 replaced by BasicMAC48_971

//BasicMAC48_649 replaced by BasicMAC48_971

//BasicMAC48_650 replaced by BasicMAC48_971

//BasicMAC48_651 replaced by BasicMAC48_971

//BasicMAC48_652 replaced by BasicMAC48_971

//BasicMAC48_653 replaced by BasicMAC48_971

//BasicMAC48_654 replaced by BasicMAC48_971

//BasicMAC48_655 replaced by BasicMAC48_971

//BasicMAC48_656 replaced by BasicMAC48_971

//BasicMAC48_657 replaced by BasicMAC48_971

//BasicMAC48_658 replaced by BasicMAC48_971

//BasicMAC48_659 replaced by BasicMAC48_971

//BasicMAC48_660 replaced by BasicMAC48_971

//BasicMAC48_661 replaced by BasicMAC48_971

//BasicMAC48_662 replaced by BasicMAC48_971

//BasicMAC48_663 replaced by BasicMAC48_971

//BasicMAC48_664 replaced by BasicMAC48_971

//BasicMAC48_665 replaced by BasicMAC48_971

//BasicMAC48_666 replaced by BasicMAC48_971

//BasicMAC48_667 replaced by BasicMAC48_971

//BasicMAC48_668 replaced by BasicMAC48_971

//BasicMAC48_669 replaced by BasicMAC48_971

//BasicMAC48_670 replaced by BasicMAC48_971

//BasicMAC48_671 replaced by BasicMAC48_971

//BasicMAC48_672 replaced by BasicMAC48_971

//BasicMAC48_673 replaced by BasicMAC48_971

//BasicMAC48_674 replaced by BasicMAC48_971

//BasicMAC48_675 replaced by BasicMAC48_971

//BasicMAC48_676 replaced by BasicMAC48_971

//BasicMAC48_677 replaced by BasicMAC48_971

//BasicMAC48_678 replaced by BasicMAC48_971

//BasicMAC48_679 replaced by BasicMAC48_971

//BasicMAC48_680 replaced by BasicMAC48_971

//BasicMAC48_681 replaced by BasicMAC48_971

//BasicMAC48_682 replaced by BasicMAC48_971

//BasicMAC48_683 replaced by BasicMAC48_971

//BasicMAC48_684 replaced by BasicMAC48_971

//BasicMAC48_685 replaced by BasicMAC48_971

//BasicMAC48_686 replaced by BasicMAC48_971

//BasicMAC48_687 replaced by BasicMAC48_971

//BasicMAC48_688 replaced by BasicMAC48_971

//BasicMAC48_689 replaced by BasicMAC48_971

//BasicMAC48_690 replaced by BasicMAC48_971

//BasicMAC48_691 replaced by BasicMAC48_971

//BasicMAC48_692 replaced by BasicMAC48_971

//BasicMAC48_693 replaced by BasicMAC48_971

//BasicMAC48_694 replaced by BasicMAC48_971

//BasicMAC48_695 replaced by BasicMAC48_971

//BasicMAC48_696 replaced by BasicMAC48_971

//BasicMAC48_697 replaced by BasicMAC48_971

//BasicMAC48_698 replaced by BasicMAC48_971

//BasicMAC48_699 replaced by BasicMAC48_971

//BasicMAC48_700 replaced by BasicMAC48_971

//BasicMAC48_701 replaced by BasicMAC48_971

//BasicMAC48_702 replaced by BasicMAC48_971

//BasicMAC48_703 replaced by BasicMAC48_971

//BasicMAC48_704 replaced by BasicMAC48_971

//BasicMAC48_705 replaced by BasicMAC48_971

//BasicMAC48_706 replaced by BasicMAC48_971

//BasicMAC48_707 replaced by BasicMAC48_971

//BasicMAC48_708 replaced by BasicMAC48_971

//BasicMAC48_709 replaced by BasicMAC48_971

//BasicMAC48_710 replaced by BasicMAC48_971

//BasicMAC48_711 replaced by BasicMAC48_971

//BasicMAC48_712 replaced by BasicMAC48_971

//BasicMAC48_713 replaced by BasicMAC48_971

//BasicMAC48_714 replaced by BasicMAC48_971

//BasicMAC48_715 replaced by BasicMAC48_971

//BasicMAC48_716 replaced by BasicMAC48_971

//BasicMAC48_717 replaced by BasicMAC48_971

//BasicMAC48_718 replaced by BasicMAC48_971

//BasicMAC48_719 replaced by BasicMAC48_971

//BasicMAC48_720 replaced by BasicMAC48_971

//BasicMAC48_721 replaced by BasicMAC48_971

//BasicMAC48_722 replaced by BasicMAC48_971

//BasicMAC48_723 replaced by BasicMAC48_971

//BasicMAC48_724 replaced by BasicMAC48_971

//BasicMAC48_725 replaced by BasicMAC48_971

//BasicMAC48_726 replaced by BasicMAC48_971

//BasicMAC48_727 replaced by BasicMAC48_971

//BasicMAC48_728 replaced by BasicMAC48_971

//BasicMAC48_729 replaced by BasicMAC48_971

//BasicMAC48_730 replaced by BasicMAC48_971

//BasicMAC48_731 replaced by BasicMAC48_971

//BasicMAC48_732 replaced by BasicMAC48_971

//BasicMAC48_733 replaced by BasicMAC48_971

//BasicMAC48_734 replaced by BasicMAC48_971

//BasicMAC48_735 replaced by BasicMAC48_971

//BasicMAC48_736 replaced by BasicMAC48_971

//BasicMAC48_737 replaced by BasicMAC48_971

//BasicMAC48_738 replaced by BasicMAC48_971

//BasicMAC48_739 replaced by BasicMAC48_971

//BasicMAC48_740 replaced by BasicMAC48_971

//BasicMAC48_741 replaced by BasicMAC48_971

//BasicMAC48_742 replaced by BasicMAC48_971

//BasicMAC48_743 replaced by BasicMAC48_971

//BasicMAC48_744 replaced by BasicMAC48_971

//BasicMAC48_745 replaced by BasicMAC48_971

//BasicMAC48_746 replaced by BasicMAC48_971

//BasicMAC48_747 replaced by BasicMAC48_971

//BasicMAC48_748 replaced by BasicMAC48_971

//BasicMAC48_749 replaced by BasicMAC48_971

//BasicMAC48_750 replaced by BasicMAC48_971

//BasicMAC48_751 replaced by BasicMAC48_971

//BasicMAC48_752 replaced by BasicMAC48_971

//BasicMAC48_753 replaced by BasicMAC48_971

//BasicMAC48_754 replaced by BasicMAC48_971

//BasicMAC48_755 replaced by BasicMAC48_971

//BasicMAC48_756 replaced by BasicMAC48_971

//BasicMAC48_757 replaced by BasicMAC48_971

//BasicMAC48_758 replaced by BasicMAC48_971

//BasicMAC48_759 replaced by BasicMAC48_971

//BasicMAC48_760 replaced by BasicMAC48_971

//BasicMAC48_761 replaced by BasicMAC48_971

//BasicMAC48_762 replaced by BasicMAC48_971

//BasicMAC48_763 replaced by BasicMAC48_971

//BasicMAC48_764 replaced by BasicMAC48_971

//BasicMAC48_765 replaced by BasicMAC48_971

//BasicMAC48_766 replaced by BasicMAC48_971

//BasicMAC48_767 replaced by BasicMAC48_971

//BasicMAC48_768 replaced by BasicMAC48_971

//BasicMAC48_769 replaced by BasicMAC48_971

//BasicMAC48_770 replaced by BasicMAC48_971

//BasicMAC48_771 replaced by BasicMAC48_971

//BasicMAC48_772 replaced by BasicMAC48_971

//BasicMAC48_773 replaced by BasicMAC48_971

//BasicMAC48_774 replaced by BasicMAC48_971

//BasicMAC48_775 replaced by BasicMAC48_971

//BasicMAC48_776 replaced by BasicMAC48_971

//BasicMAC48_777 replaced by BasicMAC48_971

//BasicMAC48_778 replaced by BasicMAC48_971

//BasicMAC48_779 replaced by BasicMAC48_971

//BasicMAC48_780 replaced by BasicMAC48_971

//BasicMAC48_781 replaced by BasicMAC48_971

//BasicMAC48_782 replaced by BasicMAC48_971

//BasicMAC48_783 replaced by BasicMAC48_971

//BasicMAC48_784 replaced by BasicMAC48_971

//BasicMAC48_785 replaced by BasicMAC48_971

//BasicMAC48_786 replaced by BasicMAC48_971

//BasicMAC48_787 replaced by BasicMAC48_971

//BasicMAC48_788 replaced by BasicMAC48_971

//BasicMAC48_789 replaced by BasicMAC48_971

//BasicMAC48_790 replaced by BasicMAC48_971

//BasicMAC48_791 replaced by BasicMAC48_971

//BasicMAC48_792 replaced by BasicMAC48_971

//BasicMAC48_793 replaced by BasicMAC48_971

//BasicMAC48_794 replaced by BasicMAC48_971

//BasicMAC48_795 replaced by BasicMAC48_971

//BasicMAC48_796 replaced by BasicMAC48_971

//BasicMAC48_797 replaced by BasicMAC48_971

//BasicMAC48_798 replaced by BasicMAC48_971

//BasicMAC48_799 replaced by BasicMAC48_971

//BasicMAC48_800 replaced by BasicMAC48_971

//BasicMAC48_801 replaced by BasicMAC48_971

//BasicMAC48_802 replaced by BasicMAC48_971

//BasicMAC48_803 replaced by BasicMAC48_971

//BasicMAC48_804 replaced by BasicMAC48_971

//BasicMAC48_805 replaced by BasicMAC48_971

//BasicMAC48_806 replaced by BasicMAC48_971

//BasicMAC48_807 replaced by BasicMAC48_971

//BasicMAC48_808 replaced by BasicMAC48_971

//BasicMAC48_809 replaced by BasicMAC48_971

//BasicMAC48_810 replaced by BasicMAC48_971

//BasicMAC48_811 replaced by BasicMAC48_971

//BasicMAC48_812 replaced by BasicMAC48_971

//BasicMAC48_813 replaced by BasicMAC48_971

//BasicMAC48_814 replaced by BasicMAC48_971

//BasicMAC48_815 replaced by BasicMAC48_971

//BasicMAC48_816 replaced by BasicMAC48_971

//BasicMAC48_817 replaced by BasicMAC48_971

//BasicMAC48_818 replaced by BasicMAC48_971

//BasicMAC48_819 replaced by BasicMAC48_971

//BasicMAC48_820 replaced by BasicMAC48_971

//BasicMAC48_821 replaced by BasicMAC48_971

//BasicMAC48_822 replaced by BasicMAC48_971

//BasicMAC48_823 replaced by BasicMAC48_971

//BasicMAC48_824 replaced by BasicMAC48_971

//BasicMAC48_825 replaced by BasicMAC48_971

//BasicMAC48_826 replaced by BasicMAC48_971

//BasicMAC48_827 replaced by BasicMAC48_971

//BasicMAC48_828 replaced by BasicMAC48_971

//BasicMAC48_829 replaced by BasicMAC48_971

//BasicMAC48_830 replaced by BasicMAC48_971

//BasicMAC48_831 replaced by BasicMAC48_971

//BasicMAC48_832 replaced by BasicMAC48_971

//BasicMAC48_833 replaced by BasicMAC48_971

//BasicMAC48_834 replaced by BasicMAC48_971

//BasicMAC48_835 replaced by BasicMAC48_971

//BasicMAC48_836 replaced by BasicMAC48_971

//BasicMAC48_837 replaced by BasicMAC48_971

//BasicMAC48_838 replaced by BasicMAC48_971

//BasicMAC48_839 replaced by BasicMAC48_971

//BasicMAC48_840 replaced by BasicMAC48_971

//BasicMAC48_841 replaced by BasicMAC48_971

//BasicMAC48_842 replaced by BasicMAC48_971

//BasicMAC48_843 replaced by BasicMAC48_971

//BasicMAC48_844 replaced by BasicMAC48_971

//BasicMAC48_845 replaced by BasicMAC48_971

//BasicMAC48_846 replaced by BasicMAC48_971

//BasicMAC48_847 replaced by BasicMAC48_971

//BasicMAC48_848 replaced by BasicMAC48_971

//BasicMAC48_849 replaced by BasicMAC48_971

//BasicMAC48_850 replaced by BasicMAC48_971

//BasicMAC48_851 replaced by BasicMAC48_971

//BasicMAC48_852 replaced by BasicMAC48_971

//BasicMAC48_853 replaced by BasicMAC48_971

//BasicMAC48_854 replaced by BasicMAC48_971

//BasicMAC48_855 replaced by BasicMAC48_971

//BasicMAC48_856 replaced by BasicMAC48_971

//BasicMAC48_857 replaced by BasicMAC48_971

//BasicMAC48_858 replaced by BasicMAC48_971

//BasicMAC48_859 replaced by BasicMAC48_971

//BasicMAC48_860 replaced by BasicMAC48_971

//BasicMAC48_861 replaced by BasicMAC48_971

//BasicMAC48_862 replaced by BasicMAC48_971

//BasicMAC48_863 replaced by BasicMAC48_971

//BasicMAC48_864 replaced by BasicMAC48_971

//BasicMAC48_865 replaced by BasicMAC48_971

//BasicMAC48_866 replaced by BasicMAC48_971

//BasicMAC48_867 replaced by BasicMAC48_971

//BasicMAC48_868 replaced by BasicMAC48_971

//BasicMAC48_869 replaced by BasicMAC48_971

//BasicMAC48_870 replaced by BasicMAC48_971

//BasicMAC48_871 replaced by BasicMAC48_971

//BasicMAC48_872 replaced by BasicMAC48_971

//BasicMAC48_873 replaced by BasicMAC48_971

//BasicMAC48_874 replaced by BasicMAC48_971

//BasicMAC48_875 replaced by BasicMAC48_971

//BasicMAC48_876 replaced by BasicMAC48_971

//BasicMAC48_877 replaced by BasicMAC48_971

//BasicMAC48_878 replaced by BasicMAC48_971

//BasicMAC48_879 replaced by BasicMAC48_971

//BasicMAC48_880 replaced by BasicMAC48_971

//BasicMAC48_881 replaced by BasicMAC48_971

//BasicMAC48_882 replaced by BasicMAC48_971

//BasicMAC48_883 replaced by BasicMAC48_971

//BasicMAC48_884 replaced by BasicMAC48_971

//BasicMAC48_885 replaced by BasicMAC48_971

//BasicMAC48_886 replaced by BasicMAC48_971

//BasicMAC48_887 replaced by BasicMAC48_971

//BasicMAC48_888 replaced by BasicMAC48_971

//BasicMAC48_889 replaced by BasicMAC48_971

//BasicMAC48_890 replaced by BasicMAC48_971

//BasicMAC48_891 replaced by BasicMAC48_971

//BasicMAC48_892 replaced by BasicMAC48_971

//BasicMAC48_893 replaced by BasicMAC48_971

//BasicMAC48_894 replaced by BasicMAC48_971

//BasicMAC48_895 replaced by BasicMAC48_971

//BasicMAC48_896 replaced by BasicMAC48_971

//BasicMAC48_897 replaced by BasicMAC48_971

//BasicMAC48_898 replaced by BasicMAC48_971

//BasicMAC48_899 replaced by BasicMAC48_971

//BasicMAC48_900 replaced by BasicMAC48_971

//BasicMAC48_901 replaced by BasicMAC48_971

//BasicMAC48_902 replaced by BasicMAC48_971

//BasicMAC48_903 replaced by BasicMAC48_971

//BasicMAC48_904 replaced by BasicMAC48_971

//BasicMAC48_905 replaced by BasicMAC48_971

//BasicMAC48_906 replaced by BasicMAC48_971

//BasicMAC48_907 replaced by BasicMAC48_971

//BasicMAC48_908 replaced by BasicMAC48_971

//BasicMAC48_909 replaced by BasicMAC48_971

//BasicMAC48_910 replaced by BasicMAC48_971

//BasicMAC48_911 replaced by BasicMAC48_971

//BasicMAC48_912 replaced by BasicMAC48_971

//BasicMAC48_913 replaced by BasicMAC48_971

//BasicMAC48_914 replaced by BasicMAC48_971

//BasicMAC48_915 replaced by BasicMAC48_971

//BasicMAC48_916 replaced by BasicMAC48_971

//BasicMAC48_917 replaced by BasicMAC48_971

//BasicMAC48_918 replaced by BasicMAC48_971

//BasicMAC48_919 replaced by BasicMAC48_971

//BasicMAC48_920 replaced by BasicMAC48_971

//BasicMAC48_921 replaced by BasicMAC48_971

//BasicMAC48_922 replaced by BasicMAC48_971

//BasicMAC48_923 replaced by BasicMAC48_971

//BasicMAC48_924 replaced by BasicMAC48_971

//BasicMAC48_925 replaced by BasicMAC48_971

//BasicMAC48_926 replaced by BasicMAC48_971

//BasicMAC48_927 replaced by BasicMAC48_971

//BasicMAC48_928 replaced by BasicMAC48_971

//BasicMAC48_929 replaced by BasicMAC48_971

//BasicMAC48_930 replaced by BasicMAC48_971

//BasicMAC48_931 replaced by BasicMAC48_971

//BasicMAC48_932 replaced by BasicMAC48_971

//BasicMAC48_933 replaced by BasicMAC48_971

//BasicMAC48_934 replaced by BasicMAC48_971

//BasicMAC48_935 replaced by BasicMAC48_971

//BasicMAC48_936 replaced by BasicMAC48_971

//BasicMAC48_937 replaced by BasicMAC48_971

//BasicMAC48_938 replaced by BasicMAC48_971

//BasicMAC48_939 replaced by BasicMAC48_971

//BasicMAC48_940 replaced by BasicMAC48_971

//BasicMAC48_941 replaced by BasicMAC48_971

//BasicMAC48_942 replaced by BasicMAC48_971

//BasicMAC48_943 replaced by BasicMAC48_971

//BasicMAC48_944 replaced by BasicMAC48_971

//BasicMAC48_945 replaced by BasicMAC48_971

//BasicMAC48_946 replaced by BasicMAC48_971

//BasicMAC48_947 replaced by BasicMAC48_971

//BasicMAC48_948 replaced by BasicMAC48_971

//BasicMAC48_949 replaced by BasicMAC48_971

//BasicMAC48_950 replaced by BasicMAC48_971

//BasicMAC48_951 replaced by BasicMAC48_971

//BasicMAC48_952 replaced by BasicMAC48_971

//BasicMAC48_953 replaced by BasicMAC48_971

//BasicMAC48_954 replaced by BasicMAC48_971

//BasicMAC48_955 replaced by BasicMAC48_971

//BasicMAC48_956 replaced by BasicMAC48_971

//BasicMAC48_957 replaced by BasicMAC48_971

//BasicMAC48_958 replaced by BasicMAC48_971

//BasicMAC48_959 replaced by BasicMAC48_971

//BasicMAC48_960 replaced by BasicMAC48_971

//BasicMAC48_961 replaced by BasicMAC48_971

//BasicMAC48_962 replaced by BasicMAC48_971

//BasicMAC48_963 replaced by BasicMAC48_971

//BasicMAC48_964 replaced by BasicMAC48_971

//BasicMAC48_965 replaced by BasicMAC48_971

//BasicMAC48_966 replaced by BasicMAC48_971

//BasicMAC48_967 replaced by BasicMAC48_971

//BasicMAC48_968 replaced by BasicMAC48_971

//BasicMAC48_969 replaced by BasicMAC48_971

//BasicMAC48_970 replaced by BasicMAC48_971

module BasicMAC48_971 (
  input      [51:0]   io_a,
  input      [50:0]   io_b,
  input      [50:0]   io_c,
  input               io_ce,
  output reg [102:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [25:0]   MACs_0_0_io_a;
  wire       [16:0]   MACs_0_0_io_b;
  reg        [16:0]   MACs_1_0_io_c;
  wire       [29:0]   MACs_0_0_io_acout;
  wire       [42:0]   MACs_0_0_io_p;
  wire       [47:0]   MACs_0_0_io_pcout;
  wire       [29:0]   MACs_0_1_io_acout;
  wire       [42:0]   MACs_0_1_io_p;
  wire       [47:0]   MACs_0_1_io_pcout;
  wire       [29:0]   MACs_0_2_io_acout;
  wire       [42:0]   MACs_0_2_io_p;
  wire       [47:0]   MACs_0_2_io_pcout;
  wire       [29:0]   MACs_1_0_io_acout;
  wire       [42:0]   MACs_1_0_io_p;
  wire       [47:0]   MACs_1_0_io_pcout;
  wire       [29:0]   MACs_1_1_io_acout;
  wire       [42:0]   MACs_1_1_io_p;
  wire       [47:0]   MACs_1_1_io_pcout;
  wire       [29:0]   MACs_1_2_io_acout;
  wire       [42:0]   MACs_1_2_io_p;
  wire       [47:0]   MACs_1_2_io_pcout;
  reg        [16:0]   _zz_io_b;
  reg        [16:0]   _zz_io_b_1;
  reg        [16:0]   _zz_io_b_2;
  reg        [16:0]   _zz_io_c;
  reg        [16:0]   _zz_io_c_1;
  reg        [16:0]   _zz_io_c_2;
  reg        [16:0]   _zz_io_c_3;
  reg        [16:0]   _zz_io_c_4;
  reg        [16:0]   _zz_io_c_5;
  reg                 _zz_io_ce;
  reg                 _zz_io_ce_1;
  reg                 _zz_io_ce_2;
  reg        [25:0]   _zz_io_a;
  reg        [25:0]   _zz_io_a_1;
  reg        [25:0]   _zz_io_a_2;
  reg        [25:0]   _zz_io_a_3;
  reg        [16:0]   _zz_io_b_3;
  reg        [16:0]   _zz_io_b_4;
  reg        [16:0]   _zz_io_b_5;
  reg        [16:0]   _zz_io_b_6;
  reg        [16:0]   _zz_io_b_7;
  reg        [16:0]   _zz_io_b_8;
  reg        [16:0]   _zz_io_b_9;
  reg        [16:0]   _zz_io_b_10;
  reg        [16:0]   _zz_io_b_11;
  reg        [16:0]   _zz_io_b_12;
  reg        [16:0]   _zz_io_b_13;
  reg        [16:0]   _zz_io_b_14;
  reg        [7:0]    _zz_io_c_6;
  reg        [16:0]   _zz_io_c_7;
  reg        [16:0]   _zz_io_c_8;
  reg        [16:0]   _zz_io_c_9;
  reg        [16:0]   _zz_io_p;
  reg        [16:0]   _zz_io_p_1;
  reg        [16:0]   _zz_io_p_2;
  reg        [16:0]   _zz_io_p_3;
  reg        [16:0]   _zz_io_p_4;
  reg        [8:0]    _zz_io_p_5;
  reg        [8:0]    _zz_io_p_6;
  reg        [8:0]    _zz_io_p_7;
  reg        [8:0]    _zz_io_p_8;
  reg        [16:0]   _zz_io_p_9;
  reg        [11:0]   _zz_io_p_10;
  reg        [6:0]    _zz_io_p_11;

  MAC_5826 MACs_0_0 (
    .io_a     (MACs_0_0_io_a[25:0]    ), //i
    .io_acin  (30'h0                  ), //i
    .io_acout (MACs_0_0_io_acout[29:0]), //o
    .io_b     (MACs_0_0_io_b[16:0]    ), //i
    .io_c     (_zz_io_c[16:0]         ), //i
    .io_ce    (_zz_io_ce              ), //i
    .io_pcin  (48'h0                  ), //i
    .io_p     (MACs_0_0_io_p[42:0]    ), //o
    .io_pcout (MACs_0_0_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_5827 MACs_0_1 (
    .io_a     (26'h0                  ), //i
    .io_acin  (MACs_0_0_io_acout[29:0]), //i
    .io_acout (MACs_0_1_io_acout[29:0]), //o
    .io_b     (_zz_io_b[16:0]         ), //i
    .io_c     (_zz_io_c_2[16:0]       ), //i
    .io_ce    (_zz_io_ce_1            ), //i
    .io_pcin  (MACs_0_0_io_pcout[47:0]), //i
    .io_p     (MACs_0_1_io_p[42:0]    ), //o
    .io_pcout (MACs_0_1_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_5827 MACs_0_2 (
    .io_a     (26'h0                  ), //i
    .io_acin  (MACs_0_1_io_acout[29:0]), //i
    .io_acout (MACs_0_2_io_acout[29:0]), //o
    .io_b     (_zz_io_b_2[16:0]       ), //i
    .io_c     (_zz_io_c_5[16:0]       ), //i
    .io_ce    (_zz_io_ce_2            ), //i
    .io_pcin  (MACs_0_1_io_pcout[47:0]), //i
    .io_p     (MACs_0_2_io_p[42:0]    ), //o
    .io_pcout (MACs_0_2_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_5826 MACs_1_0 (
    .io_a     (_zz_io_a_3[25:0]       ), //i
    .io_acin  (30'h0                  ), //i
    .io_acout (MACs_1_0_io_acout[29:0]), //o
    .io_b     (_zz_io_b_12[16:0]      ), //i
    .io_c     (MACs_1_0_io_c[16:0]    ), //i
    .io_ce    (1'b1                   ), //i
    .io_pcin  (48'h0                  ), //i
    .io_p     (MACs_1_0_io_p[42:0]    ), //o
    .io_pcout (MACs_1_0_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_5827 MACs_1_1 (
    .io_a     (26'h0                  ), //i
    .io_acin  (MACs_1_0_io_acout[29:0]), //i
    .io_acout (MACs_1_1_io_acout[29:0]), //o
    .io_b     (_zz_io_b_13[16:0]      ), //i
    .io_c     (_zz_io_c_7[16:0]       ), //i
    .io_ce    (1'b1                   ), //i
    .io_pcin  (MACs_1_0_io_pcout[47:0]), //i
    .io_p     (MACs_1_1_io_p[42:0]    ), //o
    .io_pcout (MACs_1_1_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_5827 MACs_1_2 (
    .io_a     (26'h0                  ), //i
    .io_acin  (MACs_1_1_io_acout[29:0]), //i
    .io_acout (MACs_1_2_io_acout[29:0]), //o
    .io_b     (_zz_io_b_14[16:0]      ), //i
    .io_c     (_zz_io_c_9[16:0]       ), //i
    .io_ce    (1'b1                   ), //i
    .io_pcin  (MACs_1_1_io_pcout[47:0]), //i
    .io_p     (MACs_1_2_io_p[42:0]    ), //o
    .io_pcout (MACs_1_2_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  assign MACs_0_0_io_a = io_a[25:0];
  assign MACs_0_0_io_b = io_b[16 : 0];
  always @(*) begin
    MACs_1_0_io_c[7 : 0] = _zz_io_c_6;
    MACs_1_0_io_c[16 : 8] = MACs_0_2_io_p[8 : 0];
  end

  always @(*) begin
    io_p[16 : 0] = _zz_io_p_4;
    io_p[25 : 17] = _zz_io_p_8;
    io_p[42 : 26] = _zz_io_p_9;
    io_p[47 : 43] = MACs_1_1_io_p[4 : 0];
    io_p[59 : 48] = _zz_io_p_10;
    io_p[95 : 60] = MACs_1_2_io_p[35 : 0];
    io_p[102 : 96] = _zz_io_p_11;
  end

  always @(posedge clk) begin
    _zz_io_b <= io_b[33 : 17];
    _zz_io_b_1 <= io_b[50 : 34];
    _zz_io_b_2 <= _zz_io_b_1;
    _zz_io_c <= io_c[16 : 0];
    _zz_io_c_1 <= io_c[33 : 17];
    _zz_io_c_2 <= _zz_io_c_1;
    _zz_io_c_3 <= io_c[50 : 34];
    _zz_io_c_4 <= _zz_io_c_3;
    _zz_io_c_5 <= _zz_io_c_4;
    _zz_io_ce <= io_ce;
    _zz_io_ce_1 <= _zz_io_ce;
    _zz_io_ce_2 <= _zz_io_ce_1;
    _zz_io_a <= (io_a >>> 26);
    _zz_io_a_1 <= _zz_io_a;
    _zz_io_a_2 <= _zz_io_a_1;
    _zz_io_a_3 <= _zz_io_a_2;
    _zz_io_b_3 <= MACs_0_0_io_b;
    _zz_io_b_4 <= _zz_io_b;
    _zz_io_b_5 <= _zz_io_b_2;
    _zz_io_b_6 <= _zz_io_b_3;
    _zz_io_b_7 <= _zz_io_b_4;
    _zz_io_b_8 <= _zz_io_b_5;
    _zz_io_b_9 <= _zz_io_b_6;
    _zz_io_b_10 <= _zz_io_b_7;
    _zz_io_b_11 <= _zz_io_b_8;
    _zz_io_b_12 <= _zz_io_b_9;
    _zz_io_b_13 <= _zz_io_b_10;
    _zz_io_b_14 <= _zz_io_b_11;
    _zz_io_c_6 <= MACs_0_1_io_p[16 : 9];
    _zz_io_c_7 <= MACs_0_2_io_p[25 : 9];
    _zz_io_c_8 <= MACs_0_2_io_p[42 : 26];
    _zz_io_c_9 <= _zz_io_c_8;
    _zz_io_p <= MACs_0_0_io_p[16 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= _zz_io_p_2;
    _zz_io_p_4 <= _zz_io_p_3;
    _zz_io_p_5 <= MACs_0_1_io_p[8 : 0];
    _zz_io_p_6 <= _zz_io_p_5;
    _zz_io_p_7 <= _zz_io_p_6;
    _zz_io_p_8 <= _zz_io_p_7;
    _zz_io_p_9 <= MACs_1_0_io_p[16 : 0];
    _zz_io_p_10 <= MACs_1_1_io_p[16 : 5];
    _zz_io_p_11 <= MACs_1_2_io_p[42 : 36];
  end


endmodule

//MAC_5 replaced by MAC_5827

//MAC_4 replaced by MAC_5827

//MAC_3 replaced by MAC_5826

//MAC_2 replaced by MAC_5827

//MAC_1 replaced by MAC_5827

//MAC replaced by MAC_5826

//MAC_11 replaced by MAC_5827

//MAC_10 replaced by MAC_5827

//MAC_9 replaced by MAC_5826

//MAC_8 replaced by MAC_5827

//MAC_7 replaced by MAC_5827

//MAC_6 replaced by MAC_5826

//MAC_17 replaced by MAC_5827

//MAC_16 replaced by MAC_5827

//MAC_15 replaced by MAC_5826

//MAC_14 replaced by MAC_5827

//MAC_13 replaced by MAC_5827

//MAC_12 replaced by MAC_5826

//MAC_23 replaced by MAC_5827

//MAC_22 replaced by MAC_5827

//MAC_21 replaced by MAC_5826

//MAC_20 replaced by MAC_5827

//MAC_19 replaced by MAC_5827

//MAC_18 replaced by MAC_5826

//MAC_29 replaced by MAC_5827

//MAC_28 replaced by MAC_5827

//MAC_27 replaced by MAC_5826

//MAC_26 replaced by MAC_5827

//MAC_25 replaced by MAC_5827

//MAC_24 replaced by MAC_5826

//MAC_35 replaced by MAC_5827

//MAC_34 replaced by MAC_5827

//MAC_33 replaced by MAC_5826

//MAC_32 replaced by MAC_5827

//MAC_31 replaced by MAC_5827

//MAC_30 replaced by MAC_5826

//MAC_41 replaced by MAC_5827

//MAC_40 replaced by MAC_5827

//MAC_39 replaced by MAC_5826

//MAC_38 replaced by MAC_5827

//MAC_37 replaced by MAC_5827

//MAC_36 replaced by MAC_5826

//MAC_47 replaced by MAC_5827

//MAC_46 replaced by MAC_5827

//MAC_45 replaced by MAC_5826

//MAC_44 replaced by MAC_5827

//MAC_43 replaced by MAC_5827

//MAC_42 replaced by MAC_5826

//MAC_53 replaced by MAC_5827

//MAC_52 replaced by MAC_5827

//MAC_51 replaced by MAC_5826

//MAC_50 replaced by MAC_5827

//MAC_49 replaced by MAC_5827

//MAC_48 replaced by MAC_5826

//MAC_59 replaced by MAC_5827

//MAC_58 replaced by MAC_5827

//MAC_57 replaced by MAC_5826

//MAC_56 replaced by MAC_5827

//MAC_55 replaced by MAC_5827

//MAC_54 replaced by MAC_5826

//MAC_65 replaced by MAC_5827

//MAC_64 replaced by MAC_5827

//MAC_63 replaced by MAC_5826

//MAC_62 replaced by MAC_5827

//MAC_61 replaced by MAC_5827

//MAC_60 replaced by MAC_5826

//MAC_71 replaced by MAC_5827

//MAC_70 replaced by MAC_5827

//MAC_69 replaced by MAC_5826

//MAC_68 replaced by MAC_5827

//MAC_67 replaced by MAC_5827

//MAC_66 replaced by MAC_5826

//MAC_77 replaced by MAC_5827

//MAC_76 replaced by MAC_5827

//MAC_75 replaced by MAC_5826

//MAC_74 replaced by MAC_5827

//MAC_73 replaced by MAC_5827

//MAC_72 replaced by MAC_5826

//MAC_83 replaced by MAC_5827

//MAC_82 replaced by MAC_5827

//MAC_81 replaced by MAC_5826

//MAC_80 replaced by MAC_5827

//MAC_79 replaced by MAC_5827

//MAC_78 replaced by MAC_5826

//MAC_89 replaced by MAC_5827

//MAC_88 replaced by MAC_5827

//MAC_87 replaced by MAC_5826

//MAC_86 replaced by MAC_5827

//MAC_85 replaced by MAC_5827

//MAC_84 replaced by MAC_5826

//MAC_95 replaced by MAC_5827

//MAC_94 replaced by MAC_5827

//MAC_93 replaced by MAC_5826

//MAC_92 replaced by MAC_5827

//MAC_91 replaced by MAC_5827

//MAC_90 replaced by MAC_5826

//MAC_101 replaced by MAC_5827

//MAC_100 replaced by MAC_5827

//MAC_99 replaced by MAC_5826

//MAC_98 replaced by MAC_5827

//MAC_97 replaced by MAC_5827

//MAC_96 replaced by MAC_5826

//MAC_107 replaced by MAC_5827

//MAC_106 replaced by MAC_5827

//MAC_105 replaced by MAC_5826

//MAC_104 replaced by MAC_5827

//MAC_103 replaced by MAC_5827

//MAC_102 replaced by MAC_5826

//MAC_113 replaced by MAC_5827

//MAC_112 replaced by MAC_5827

//MAC_111 replaced by MAC_5826

//MAC_110 replaced by MAC_5827

//MAC_109 replaced by MAC_5827

//MAC_108 replaced by MAC_5826

//MAC_119 replaced by MAC_5827

//MAC_118 replaced by MAC_5827

//MAC_117 replaced by MAC_5826

//MAC_116 replaced by MAC_5827

//MAC_115 replaced by MAC_5827

//MAC_114 replaced by MAC_5826

//MAC_125 replaced by MAC_5827

//MAC_124 replaced by MAC_5827

//MAC_123 replaced by MAC_5826

//MAC_122 replaced by MAC_5827

//MAC_121 replaced by MAC_5827

//MAC_120 replaced by MAC_5826

//MAC_131 replaced by MAC_5827

//MAC_130 replaced by MAC_5827

//MAC_129 replaced by MAC_5826

//MAC_128 replaced by MAC_5827

//MAC_127 replaced by MAC_5827

//MAC_126 replaced by MAC_5826

//MAC_137 replaced by MAC_5827

//MAC_136 replaced by MAC_5827

//MAC_135 replaced by MAC_5826

//MAC_134 replaced by MAC_5827

//MAC_133 replaced by MAC_5827

//MAC_132 replaced by MAC_5826

//MAC_143 replaced by MAC_5827

//MAC_142 replaced by MAC_5827

//MAC_141 replaced by MAC_5826

//MAC_140 replaced by MAC_5827

//MAC_139 replaced by MAC_5827

//MAC_138 replaced by MAC_5826

//MAC_149 replaced by MAC_5827

//MAC_148 replaced by MAC_5827

//MAC_147 replaced by MAC_5826

//MAC_146 replaced by MAC_5827

//MAC_145 replaced by MAC_5827

//MAC_144 replaced by MAC_5826

//MAC_155 replaced by MAC_5827

//MAC_154 replaced by MAC_5827

//MAC_153 replaced by MAC_5826

//MAC_152 replaced by MAC_5827

//MAC_151 replaced by MAC_5827

//MAC_150 replaced by MAC_5826

//MAC_161 replaced by MAC_5827

//MAC_160 replaced by MAC_5827

//MAC_159 replaced by MAC_5826

//MAC_158 replaced by MAC_5827

//MAC_157 replaced by MAC_5827

//MAC_156 replaced by MAC_5826

//MAC_167 replaced by MAC_5827

//MAC_166 replaced by MAC_5827

//MAC_165 replaced by MAC_5826

//MAC_164 replaced by MAC_5827

//MAC_163 replaced by MAC_5827

//MAC_162 replaced by MAC_5826

//MAC_173 replaced by MAC_5827

//MAC_172 replaced by MAC_5827

//MAC_171 replaced by MAC_5826

//MAC_170 replaced by MAC_5827

//MAC_169 replaced by MAC_5827

//MAC_168 replaced by MAC_5826

//MAC_179 replaced by MAC_5827

//MAC_178 replaced by MAC_5827

//MAC_177 replaced by MAC_5826

//MAC_176 replaced by MAC_5827

//MAC_175 replaced by MAC_5827

//MAC_174 replaced by MAC_5826

//MAC_185 replaced by MAC_5827

//MAC_184 replaced by MAC_5827

//MAC_183 replaced by MAC_5826

//MAC_182 replaced by MAC_5827

//MAC_181 replaced by MAC_5827

//MAC_180 replaced by MAC_5826

//MAC_191 replaced by MAC_5827

//MAC_190 replaced by MAC_5827

//MAC_189 replaced by MAC_5826

//MAC_188 replaced by MAC_5827

//MAC_187 replaced by MAC_5827

//MAC_186 replaced by MAC_5826

//MAC_197 replaced by MAC_5827

//MAC_196 replaced by MAC_5827

//MAC_195 replaced by MAC_5826

//MAC_194 replaced by MAC_5827

//MAC_193 replaced by MAC_5827

//MAC_192 replaced by MAC_5826

//MAC_203 replaced by MAC_5827

//MAC_202 replaced by MAC_5827

//MAC_201 replaced by MAC_5826

//MAC_200 replaced by MAC_5827

//MAC_199 replaced by MAC_5827

//MAC_198 replaced by MAC_5826

//MAC_209 replaced by MAC_5827

//MAC_208 replaced by MAC_5827

//MAC_207 replaced by MAC_5826

//MAC_206 replaced by MAC_5827

//MAC_205 replaced by MAC_5827

//MAC_204 replaced by MAC_5826

//MAC_215 replaced by MAC_5827

//MAC_214 replaced by MAC_5827

//MAC_213 replaced by MAC_5826

//MAC_212 replaced by MAC_5827

//MAC_211 replaced by MAC_5827

//MAC_210 replaced by MAC_5826

//MAC_221 replaced by MAC_5827

//MAC_220 replaced by MAC_5827

//MAC_219 replaced by MAC_5826

//MAC_218 replaced by MAC_5827

//MAC_217 replaced by MAC_5827

//MAC_216 replaced by MAC_5826

//MAC_227 replaced by MAC_5827

//MAC_226 replaced by MAC_5827

//MAC_225 replaced by MAC_5826

//MAC_224 replaced by MAC_5827

//MAC_223 replaced by MAC_5827

//MAC_222 replaced by MAC_5826

//MAC_233 replaced by MAC_5827

//MAC_232 replaced by MAC_5827

//MAC_231 replaced by MAC_5826

//MAC_230 replaced by MAC_5827

//MAC_229 replaced by MAC_5827

//MAC_228 replaced by MAC_5826

//MAC_239 replaced by MAC_5827

//MAC_238 replaced by MAC_5827

//MAC_237 replaced by MAC_5826

//MAC_236 replaced by MAC_5827

//MAC_235 replaced by MAC_5827

//MAC_234 replaced by MAC_5826

//MAC_245 replaced by MAC_5827

//MAC_244 replaced by MAC_5827

//MAC_243 replaced by MAC_5826

//MAC_242 replaced by MAC_5827

//MAC_241 replaced by MAC_5827

//MAC_240 replaced by MAC_5826

//MAC_251 replaced by MAC_5827

//MAC_250 replaced by MAC_5827

//MAC_249 replaced by MAC_5826

//MAC_248 replaced by MAC_5827

//MAC_247 replaced by MAC_5827

//MAC_246 replaced by MAC_5826

//MAC_257 replaced by MAC_5827

//MAC_256 replaced by MAC_5827

//MAC_255 replaced by MAC_5826

//MAC_254 replaced by MAC_5827

//MAC_253 replaced by MAC_5827

//MAC_252 replaced by MAC_5826

//MAC_263 replaced by MAC_5827

//MAC_262 replaced by MAC_5827

//MAC_261 replaced by MAC_5826

//MAC_260 replaced by MAC_5827

//MAC_259 replaced by MAC_5827

//MAC_258 replaced by MAC_5826

//MAC_269 replaced by MAC_5827

//MAC_268 replaced by MAC_5827

//MAC_267 replaced by MAC_5826

//MAC_266 replaced by MAC_5827

//MAC_265 replaced by MAC_5827

//MAC_264 replaced by MAC_5826

//MAC_275 replaced by MAC_5827

//MAC_274 replaced by MAC_5827

//MAC_273 replaced by MAC_5826

//MAC_272 replaced by MAC_5827

//MAC_271 replaced by MAC_5827

//MAC_270 replaced by MAC_5826

//MAC_281 replaced by MAC_5827

//MAC_280 replaced by MAC_5827

//MAC_279 replaced by MAC_5826

//MAC_278 replaced by MAC_5827

//MAC_277 replaced by MAC_5827

//MAC_276 replaced by MAC_5826

//MAC_287 replaced by MAC_5827

//MAC_286 replaced by MAC_5827

//MAC_285 replaced by MAC_5826

//MAC_284 replaced by MAC_5827

//MAC_283 replaced by MAC_5827

//MAC_282 replaced by MAC_5826

//MAC_293 replaced by MAC_5827

//MAC_292 replaced by MAC_5827

//MAC_291 replaced by MAC_5826

//MAC_290 replaced by MAC_5827

//MAC_289 replaced by MAC_5827

//MAC_288 replaced by MAC_5826

//MAC_299 replaced by MAC_5827

//MAC_298 replaced by MAC_5827

//MAC_297 replaced by MAC_5826

//MAC_296 replaced by MAC_5827

//MAC_295 replaced by MAC_5827

//MAC_294 replaced by MAC_5826

//MAC_305 replaced by MAC_5827

//MAC_304 replaced by MAC_5827

//MAC_303 replaced by MAC_5826

//MAC_302 replaced by MAC_5827

//MAC_301 replaced by MAC_5827

//MAC_300 replaced by MAC_5826

//MAC_311 replaced by MAC_5827

//MAC_310 replaced by MAC_5827

//MAC_309 replaced by MAC_5826

//MAC_308 replaced by MAC_5827

//MAC_307 replaced by MAC_5827

//MAC_306 replaced by MAC_5826

//MAC_317 replaced by MAC_5827

//MAC_316 replaced by MAC_5827

//MAC_315 replaced by MAC_5826

//MAC_314 replaced by MAC_5827

//MAC_313 replaced by MAC_5827

//MAC_312 replaced by MAC_5826

//MAC_323 replaced by MAC_5827

//MAC_322 replaced by MAC_5827

//MAC_321 replaced by MAC_5826

//MAC_320 replaced by MAC_5827

//MAC_319 replaced by MAC_5827

//MAC_318 replaced by MAC_5826

//MAC_329 replaced by MAC_5827

//MAC_328 replaced by MAC_5827

//MAC_327 replaced by MAC_5826

//MAC_326 replaced by MAC_5827

//MAC_325 replaced by MAC_5827

//MAC_324 replaced by MAC_5826

//MAC_335 replaced by MAC_5827

//MAC_334 replaced by MAC_5827

//MAC_333 replaced by MAC_5826

//MAC_332 replaced by MAC_5827

//MAC_331 replaced by MAC_5827

//MAC_330 replaced by MAC_5826

//MAC_341 replaced by MAC_5827

//MAC_340 replaced by MAC_5827

//MAC_339 replaced by MAC_5826

//MAC_338 replaced by MAC_5827

//MAC_337 replaced by MAC_5827

//MAC_336 replaced by MAC_5826

//MAC_347 replaced by MAC_5827

//MAC_346 replaced by MAC_5827

//MAC_345 replaced by MAC_5826

//MAC_344 replaced by MAC_5827

//MAC_343 replaced by MAC_5827

//MAC_342 replaced by MAC_5826

//MAC_353 replaced by MAC_5827

//MAC_352 replaced by MAC_5827

//MAC_351 replaced by MAC_5826

//MAC_350 replaced by MAC_5827

//MAC_349 replaced by MAC_5827

//MAC_348 replaced by MAC_5826

//MAC_359 replaced by MAC_5827

//MAC_358 replaced by MAC_5827

//MAC_357 replaced by MAC_5826

//MAC_356 replaced by MAC_5827

//MAC_355 replaced by MAC_5827

//MAC_354 replaced by MAC_5826

//MAC_365 replaced by MAC_5827

//MAC_364 replaced by MAC_5827

//MAC_363 replaced by MAC_5826

//MAC_362 replaced by MAC_5827

//MAC_361 replaced by MAC_5827

//MAC_360 replaced by MAC_5826

//MAC_371 replaced by MAC_5827

//MAC_370 replaced by MAC_5827

//MAC_369 replaced by MAC_5826

//MAC_368 replaced by MAC_5827

//MAC_367 replaced by MAC_5827

//MAC_366 replaced by MAC_5826

//MAC_377 replaced by MAC_5827

//MAC_376 replaced by MAC_5827

//MAC_375 replaced by MAC_5826

//MAC_374 replaced by MAC_5827

//MAC_373 replaced by MAC_5827

//MAC_372 replaced by MAC_5826

//MAC_383 replaced by MAC_5827

//MAC_382 replaced by MAC_5827

//MAC_381 replaced by MAC_5826

//MAC_380 replaced by MAC_5827

//MAC_379 replaced by MAC_5827

//MAC_378 replaced by MAC_5826

//MAC_389 replaced by MAC_5827

//MAC_388 replaced by MAC_5827

//MAC_387 replaced by MAC_5826

//MAC_386 replaced by MAC_5827

//MAC_385 replaced by MAC_5827

//MAC_384 replaced by MAC_5826

//MAC_395 replaced by MAC_5827

//MAC_394 replaced by MAC_5827

//MAC_393 replaced by MAC_5826

//MAC_392 replaced by MAC_5827

//MAC_391 replaced by MAC_5827

//MAC_390 replaced by MAC_5826

//MAC_401 replaced by MAC_5827

//MAC_400 replaced by MAC_5827

//MAC_399 replaced by MAC_5826

//MAC_398 replaced by MAC_5827

//MAC_397 replaced by MAC_5827

//MAC_396 replaced by MAC_5826

//MAC_407 replaced by MAC_5827

//MAC_406 replaced by MAC_5827

//MAC_405 replaced by MAC_5826

//MAC_404 replaced by MAC_5827

//MAC_403 replaced by MAC_5827

//MAC_402 replaced by MAC_5826

//MAC_413 replaced by MAC_5827

//MAC_412 replaced by MAC_5827

//MAC_411 replaced by MAC_5826

//MAC_410 replaced by MAC_5827

//MAC_409 replaced by MAC_5827

//MAC_408 replaced by MAC_5826

//MAC_419 replaced by MAC_5827

//MAC_418 replaced by MAC_5827

//MAC_417 replaced by MAC_5826

//MAC_416 replaced by MAC_5827

//MAC_415 replaced by MAC_5827

//MAC_414 replaced by MAC_5826

//MAC_425 replaced by MAC_5827

//MAC_424 replaced by MAC_5827

//MAC_423 replaced by MAC_5826

//MAC_422 replaced by MAC_5827

//MAC_421 replaced by MAC_5827

//MAC_420 replaced by MAC_5826

//MAC_431 replaced by MAC_5827

//MAC_430 replaced by MAC_5827

//MAC_429 replaced by MAC_5826

//MAC_428 replaced by MAC_5827

//MAC_427 replaced by MAC_5827

//MAC_426 replaced by MAC_5826

//MAC_437 replaced by MAC_5827

//MAC_436 replaced by MAC_5827

//MAC_435 replaced by MAC_5826

//MAC_434 replaced by MAC_5827

//MAC_433 replaced by MAC_5827

//MAC_432 replaced by MAC_5826

//MAC_443 replaced by MAC_5827

//MAC_442 replaced by MAC_5827

//MAC_441 replaced by MAC_5826

//MAC_440 replaced by MAC_5827

//MAC_439 replaced by MAC_5827

//MAC_438 replaced by MAC_5826

//MAC_449 replaced by MAC_5827

//MAC_448 replaced by MAC_5827

//MAC_447 replaced by MAC_5826

//MAC_446 replaced by MAC_5827

//MAC_445 replaced by MAC_5827

//MAC_444 replaced by MAC_5826

//MAC_455 replaced by MAC_5827

//MAC_454 replaced by MAC_5827

//MAC_453 replaced by MAC_5826

//MAC_452 replaced by MAC_5827

//MAC_451 replaced by MAC_5827

//MAC_450 replaced by MAC_5826

//MAC_461 replaced by MAC_5827

//MAC_460 replaced by MAC_5827

//MAC_459 replaced by MAC_5826

//MAC_458 replaced by MAC_5827

//MAC_457 replaced by MAC_5827

//MAC_456 replaced by MAC_5826

//MAC_467 replaced by MAC_5827

//MAC_466 replaced by MAC_5827

//MAC_465 replaced by MAC_5826

//MAC_464 replaced by MAC_5827

//MAC_463 replaced by MAC_5827

//MAC_462 replaced by MAC_5826

//MAC_473 replaced by MAC_5827

//MAC_472 replaced by MAC_5827

//MAC_471 replaced by MAC_5826

//MAC_470 replaced by MAC_5827

//MAC_469 replaced by MAC_5827

//MAC_468 replaced by MAC_5826

//MAC_479 replaced by MAC_5827

//MAC_478 replaced by MAC_5827

//MAC_477 replaced by MAC_5826

//MAC_476 replaced by MAC_5827

//MAC_475 replaced by MAC_5827

//MAC_474 replaced by MAC_5826

//MAC_485 replaced by MAC_5827

//MAC_484 replaced by MAC_5827

//MAC_483 replaced by MAC_5826

//MAC_482 replaced by MAC_5827

//MAC_481 replaced by MAC_5827

//MAC_480 replaced by MAC_5826

//MAC_491 replaced by MAC_5827

//MAC_490 replaced by MAC_5827

//MAC_489 replaced by MAC_5826

//MAC_488 replaced by MAC_5827

//MAC_487 replaced by MAC_5827

//MAC_486 replaced by MAC_5826

//MAC_497 replaced by MAC_5827

//MAC_496 replaced by MAC_5827

//MAC_495 replaced by MAC_5826

//MAC_494 replaced by MAC_5827

//MAC_493 replaced by MAC_5827

//MAC_492 replaced by MAC_5826

//MAC_503 replaced by MAC_5827

//MAC_502 replaced by MAC_5827

//MAC_501 replaced by MAC_5826

//MAC_500 replaced by MAC_5827

//MAC_499 replaced by MAC_5827

//MAC_498 replaced by MAC_5826

//MAC_509 replaced by MAC_5827

//MAC_508 replaced by MAC_5827

//MAC_507 replaced by MAC_5826

//MAC_506 replaced by MAC_5827

//MAC_505 replaced by MAC_5827

//MAC_504 replaced by MAC_5826

//MAC_515 replaced by MAC_5827

//MAC_514 replaced by MAC_5827

//MAC_513 replaced by MAC_5826

//MAC_512 replaced by MAC_5827

//MAC_511 replaced by MAC_5827

//MAC_510 replaced by MAC_5826

//MAC_521 replaced by MAC_5827

//MAC_520 replaced by MAC_5827

//MAC_519 replaced by MAC_5826

//MAC_518 replaced by MAC_5827

//MAC_517 replaced by MAC_5827

//MAC_516 replaced by MAC_5826

//MAC_527 replaced by MAC_5827

//MAC_526 replaced by MAC_5827

//MAC_525 replaced by MAC_5826

//MAC_524 replaced by MAC_5827

//MAC_523 replaced by MAC_5827

//MAC_522 replaced by MAC_5826

//MAC_533 replaced by MAC_5827

//MAC_532 replaced by MAC_5827

//MAC_531 replaced by MAC_5826

//MAC_530 replaced by MAC_5827

//MAC_529 replaced by MAC_5827

//MAC_528 replaced by MAC_5826

//MAC_539 replaced by MAC_5827

//MAC_538 replaced by MAC_5827

//MAC_537 replaced by MAC_5826

//MAC_536 replaced by MAC_5827

//MAC_535 replaced by MAC_5827

//MAC_534 replaced by MAC_5826

//MAC_545 replaced by MAC_5827

//MAC_544 replaced by MAC_5827

//MAC_543 replaced by MAC_5826

//MAC_542 replaced by MAC_5827

//MAC_541 replaced by MAC_5827

//MAC_540 replaced by MAC_5826

//MAC_551 replaced by MAC_5827

//MAC_550 replaced by MAC_5827

//MAC_549 replaced by MAC_5826

//MAC_548 replaced by MAC_5827

//MAC_547 replaced by MAC_5827

//MAC_546 replaced by MAC_5826

//MAC_557 replaced by MAC_5827

//MAC_556 replaced by MAC_5827

//MAC_555 replaced by MAC_5826

//MAC_554 replaced by MAC_5827

//MAC_553 replaced by MAC_5827

//MAC_552 replaced by MAC_5826

//MAC_563 replaced by MAC_5827

//MAC_562 replaced by MAC_5827

//MAC_561 replaced by MAC_5826

//MAC_560 replaced by MAC_5827

//MAC_559 replaced by MAC_5827

//MAC_558 replaced by MAC_5826

//MAC_569 replaced by MAC_5827

//MAC_568 replaced by MAC_5827

//MAC_567 replaced by MAC_5826

//MAC_566 replaced by MAC_5827

//MAC_565 replaced by MAC_5827

//MAC_564 replaced by MAC_5826

//MAC_575 replaced by MAC_5827

//MAC_574 replaced by MAC_5827

//MAC_573 replaced by MAC_5826

//MAC_572 replaced by MAC_5827

//MAC_571 replaced by MAC_5827

//MAC_570 replaced by MAC_5826

//MAC_581 replaced by MAC_5827

//MAC_580 replaced by MAC_5827

//MAC_579 replaced by MAC_5826

//MAC_578 replaced by MAC_5827

//MAC_577 replaced by MAC_5827

//MAC_576 replaced by MAC_5826

//MAC_587 replaced by MAC_5827

//MAC_586 replaced by MAC_5827

//MAC_585 replaced by MAC_5826

//MAC_584 replaced by MAC_5827

//MAC_583 replaced by MAC_5827

//MAC_582 replaced by MAC_5826

//MAC_593 replaced by MAC_5827

//MAC_592 replaced by MAC_5827

//MAC_591 replaced by MAC_5826

//MAC_590 replaced by MAC_5827

//MAC_589 replaced by MAC_5827

//MAC_588 replaced by MAC_5826

//MAC_599 replaced by MAC_5827

//MAC_598 replaced by MAC_5827

//MAC_597 replaced by MAC_5826

//MAC_596 replaced by MAC_5827

//MAC_595 replaced by MAC_5827

//MAC_594 replaced by MAC_5826

//MAC_605 replaced by MAC_5827

//MAC_604 replaced by MAC_5827

//MAC_603 replaced by MAC_5826

//MAC_602 replaced by MAC_5827

//MAC_601 replaced by MAC_5827

//MAC_600 replaced by MAC_5826

//MAC_611 replaced by MAC_5827

//MAC_610 replaced by MAC_5827

//MAC_609 replaced by MAC_5826

//MAC_608 replaced by MAC_5827

//MAC_607 replaced by MAC_5827

//MAC_606 replaced by MAC_5826

//MAC_617 replaced by MAC_5827

//MAC_616 replaced by MAC_5827

//MAC_615 replaced by MAC_5826

//MAC_614 replaced by MAC_5827

//MAC_613 replaced by MAC_5827

//MAC_612 replaced by MAC_5826

//MAC_623 replaced by MAC_5827

//MAC_622 replaced by MAC_5827

//MAC_621 replaced by MAC_5826

//MAC_620 replaced by MAC_5827

//MAC_619 replaced by MAC_5827

//MAC_618 replaced by MAC_5826

//MAC_629 replaced by MAC_5827

//MAC_628 replaced by MAC_5827

//MAC_627 replaced by MAC_5826

//MAC_626 replaced by MAC_5827

//MAC_625 replaced by MAC_5827

//MAC_624 replaced by MAC_5826

//MAC_635 replaced by MAC_5827

//MAC_634 replaced by MAC_5827

//MAC_633 replaced by MAC_5826

//MAC_632 replaced by MAC_5827

//MAC_631 replaced by MAC_5827

//MAC_630 replaced by MAC_5826

//MAC_641 replaced by MAC_5827

//MAC_640 replaced by MAC_5827

//MAC_639 replaced by MAC_5826

//MAC_638 replaced by MAC_5827

//MAC_637 replaced by MAC_5827

//MAC_636 replaced by MAC_5826

//MAC_647 replaced by MAC_5827

//MAC_646 replaced by MAC_5827

//MAC_645 replaced by MAC_5826

//MAC_644 replaced by MAC_5827

//MAC_643 replaced by MAC_5827

//MAC_642 replaced by MAC_5826

//MAC_653 replaced by MAC_5827

//MAC_652 replaced by MAC_5827

//MAC_651 replaced by MAC_5826

//MAC_650 replaced by MAC_5827

//MAC_649 replaced by MAC_5827

//MAC_648 replaced by MAC_5826

//MAC_659 replaced by MAC_5827

//MAC_658 replaced by MAC_5827

//MAC_657 replaced by MAC_5826

//MAC_656 replaced by MAC_5827

//MAC_655 replaced by MAC_5827

//MAC_654 replaced by MAC_5826

//MAC_665 replaced by MAC_5827

//MAC_664 replaced by MAC_5827

//MAC_663 replaced by MAC_5826

//MAC_662 replaced by MAC_5827

//MAC_661 replaced by MAC_5827

//MAC_660 replaced by MAC_5826

//MAC_671 replaced by MAC_5827

//MAC_670 replaced by MAC_5827

//MAC_669 replaced by MAC_5826

//MAC_668 replaced by MAC_5827

//MAC_667 replaced by MAC_5827

//MAC_666 replaced by MAC_5826

//MAC_677 replaced by MAC_5827

//MAC_676 replaced by MAC_5827

//MAC_675 replaced by MAC_5826

//MAC_674 replaced by MAC_5827

//MAC_673 replaced by MAC_5827

//MAC_672 replaced by MAC_5826

//MAC_683 replaced by MAC_5827

//MAC_682 replaced by MAC_5827

//MAC_681 replaced by MAC_5826

//MAC_680 replaced by MAC_5827

//MAC_679 replaced by MAC_5827

//MAC_678 replaced by MAC_5826

//MAC_689 replaced by MAC_5827

//MAC_688 replaced by MAC_5827

//MAC_687 replaced by MAC_5826

//MAC_686 replaced by MAC_5827

//MAC_685 replaced by MAC_5827

//MAC_684 replaced by MAC_5826

//MAC_695 replaced by MAC_5827

//MAC_694 replaced by MAC_5827

//MAC_693 replaced by MAC_5826

//MAC_692 replaced by MAC_5827

//MAC_691 replaced by MAC_5827

//MAC_690 replaced by MAC_5826

//MAC_701 replaced by MAC_5827

//MAC_700 replaced by MAC_5827

//MAC_699 replaced by MAC_5826

//MAC_698 replaced by MAC_5827

//MAC_697 replaced by MAC_5827

//MAC_696 replaced by MAC_5826

//MAC_707 replaced by MAC_5827

//MAC_706 replaced by MAC_5827

//MAC_705 replaced by MAC_5826

//MAC_704 replaced by MAC_5827

//MAC_703 replaced by MAC_5827

//MAC_702 replaced by MAC_5826

//MAC_713 replaced by MAC_5827

//MAC_712 replaced by MAC_5827

//MAC_711 replaced by MAC_5826

//MAC_710 replaced by MAC_5827

//MAC_709 replaced by MAC_5827

//MAC_708 replaced by MAC_5826

//MAC_719 replaced by MAC_5827

//MAC_718 replaced by MAC_5827

//MAC_717 replaced by MAC_5826

//MAC_716 replaced by MAC_5827

//MAC_715 replaced by MAC_5827

//MAC_714 replaced by MAC_5826

//MAC_725 replaced by MAC_5827

//MAC_724 replaced by MAC_5827

//MAC_723 replaced by MAC_5826

//MAC_722 replaced by MAC_5827

//MAC_721 replaced by MAC_5827

//MAC_720 replaced by MAC_5826

//MAC_731 replaced by MAC_5827

//MAC_730 replaced by MAC_5827

//MAC_729 replaced by MAC_5826

//MAC_728 replaced by MAC_5827

//MAC_727 replaced by MAC_5827

//MAC_726 replaced by MAC_5826

//MAC_737 replaced by MAC_5827

//MAC_736 replaced by MAC_5827

//MAC_735 replaced by MAC_5826

//MAC_734 replaced by MAC_5827

//MAC_733 replaced by MAC_5827

//MAC_732 replaced by MAC_5826

//MAC_743 replaced by MAC_5827

//MAC_742 replaced by MAC_5827

//MAC_741 replaced by MAC_5826

//MAC_740 replaced by MAC_5827

//MAC_739 replaced by MAC_5827

//MAC_738 replaced by MAC_5826

//MAC_749 replaced by MAC_5827

//MAC_748 replaced by MAC_5827

//MAC_747 replaced by MAC_5826

//MAC_746 replaced by MAC_5827

//MAC_745 replaced by MAC_5827

//MAC_744 replaced by MAC_5826

//MAC_755 replaced by MAC_5827

//MAC_754 replaced by MAC_5827

//MAC_753 replaced by MAC_5826

//MAC_752 replaced by MAC_5827

//MAC_751 replaced by MAC_5827

//MAC_750 replaced by MAC_5826

//MAC_761 replaced by MAC_5827

//MAC_760 replaced by MAC_5827

//MAC_759 replaced by MAC_5826

//MAC_758 replaced by MAC_5827

//MAC_757 replaced by MAC_5827

//MAC_756 replaced by MAC_5826

//MAC_767 replaced by MAC_5827

//MAC_766 replaced by MAC_5827

//MAC_765 replaced by MAC_5826

//MAC_764 replaced by MAC_5827

//MAC_763 replaced by MAC_5827

//MAC_762 replaced by MAC_5826

//MAC_773 replaced by MAC_5827

//MAC_772 replaced by MAC_5827

//MAC_771 replaced by MAC_5826

//MAC_770 replaced by MAC_5827

//MAC_769 replaced by MAC_5827

//MAC_768 replaced by MAC_5826

//MAC_779 replaced by MAC_5827

//MAC_778 replaced by MAC_5827

//MAC_777 replaced by MAC_5826

//MAC_776 replaced by MAC_5827

//MAC_775 replaced by MAC_5827

//MAC_774 replaced by MAC_5826

//MAC_785 replaced by MAC_5827

//MAC_784 replaced by MAC_5827

//MAC_783 replaced by MAC_5826

//MAC_782 replaced by MAC_5827

//MAC_781 replaced by MAC_5827

//MAC_780 replaced by MAC_5826

//MAC_791 replaced by MAC_5827

//MAC_790 replaced by MAC_5827

//MAC_789 replaced by MAC_5826

//MAC_788 replaced by MAC_5827

//MAC_787 replaced by MAC_5827

//MAC_786 replaced by MAC_5826

//MAC_797 replaced by MAC_5827

//MAC_796 replaced by MAC_5827

//MAC_795 replaced by MAC_5826

//MAC_794 replaced by MAC_5827

//MAC_793 replaced by MAC_5827

//MAC_792 replaced by MAC_5826

//MAC_803 replaced by MAC_5827

//MAC_802 replaced by MAC_5827

//MAC_801 replaced by MAC_5826

//MAC_800 replaced by MAC_5827

//MAC_799 replaced by MAC_5827

//MAC_798 replaced by MAC_5826

//MAC_809 replaced by MAC_5827

//MAC_808 replaced by MAC_5827

//MAC_807 replaced by MAC_5826

//MAC_806 replaced by MAC_5827

//MAC_805 replaced by MAC_5827

//MAC_804 replaced by MAC_5826

//MAC_815 replaced by MAC_5827

//MAC_814 replaced by MAC_5827

//MAC_813 replaced by MAC_5826

//MAC_812 replaced by MAC_5827

//MAC_811 replaced by MAC_5827

//MAC_810 replaced by MAC_5826

//MAC_821 replaced by MAC_5827

//MAC_820 replaced by MAC_5827

//MAC_819 replaced by MAC_5826

//MAC_818 replaced by MAC_5827

//MAC_817 replaced by MAC_5827

//MAC_816 replaced by MAC_5826

//MAC_827 replaced by MAC_5827

//MAC_826 replaced by MAC_5827

//MAC_825 replaced by MAC_5826

//MAC_824 replaced by MAC_5827

//MAC_823 replaced by MAC_5827

//MAC_822 replaced by MAC_5826

//MAC_833 replaced by MAC_5827

//MAC_832 replaced by MAC_5827

//MAC_831 replaced by MAC_5826

//MAC_830 replaced by MAC_5827

//MAC_829 replaced by MAC_5827

//MAC_828 replaced by MAC_5826

//MAC_839 replaced by MAC_5827

//MAC_838 replaced by MAC_5827

//MAC_837 replaced by MAC_5826

//MAC_836 replaced by MAC_5827

//MAC_835 replaced by MAC_5827

//MAC_834 replaced by MAC_5826

//MAC_845 replaced by MAC_5827

//MAC_844 replaced by MAC_5827

//MAC_843 replaced by MAC_5826

//MAC_842 replaced by MAC_5827

//MAC_841 replaced by MAC_5827

//MAC_840 replaced by MAC_5826

//MAC_851 replaced by MAC_5827

//MAC_850 replaced by MAC_5827

//MAC_849 replaced by MAC_5826

//MAC_848 replaced by MAC_5827

//MAC_847 replaced by MAC_5827

//MAC_846 replaced by MAC_5826

//MAC_857 replaced by MAC_5827

//MAC_856 replaced by MAC_5827

//MAC_855 replaced by MAC_5826

//MAC_854 replaced by MAC_5827

//MAC_853 replaced by MAC_5827

//MAC_852 replaced by MAC_5826

//MAC_863 replaced by MAC_5827

//MAC_862 replaced by MAC_5827

//MAC_861 replaced by MAC_5826

//MAC_860 replaced by MAC_5827

//MAC_859 replaced by MAC_5827

//MAC_858 replaced by MAC_5826

//MAC_869 replaced by MAC_5827

//MAC_868 replaced by MAC_5827

//MAC_867 replaced by MAC_5826

//MAC_866 replaced by MAC_5827

//MAC_865 replaced by MAC_5827

//MAC_864 replaced by MAC_5826

//MAC_875 replaced by MAC_5827

//MAC_874 replaced by MAC_5827

//MAC_873 replaced by MAC_5826

//MAC_872 replaced by MAC_5827

//MAC_871 replaced by MAC_5827

//MAC_870 replaced by MAC_5826

//MAC_881 replaced by MAC_5827

//MAC_880 replaced by MAC_5827

//MAC_879 replaced by MAC_5826

//MAC_878 replaced by MAC_5827

//MAC_877 replaced by MAC_5827

//MAC_876 replaced by MAC_5826

//MAC_887 replaced by MAC_5827

//MAC_886 replaced by MAC_5827

//MAC_885 replaced by MAC_5826

//MAC_884 replaced by MAC_5827

//MAC_883 replaced by MAC_5827

//MAC_882 replaced by MAC_5826

//MAC_893 replaced by MAC_5827

//MAC_892 replaced by MAC_5827

//MAC_891 replaced by MAC_5826

//MAC_890 replaced by MAC_5827

//MAC_889 replaced by MAC_5827

//MAC_888 replaced by MAC_5826

//MAC_899 replaced by MAC_5827

//MAC_898 replaced by MAC_5827

//MAC_897 replaced by MAC_5826

//MAC_896 replaced by MAC_5827

//MAC_895 replaced by MAC_5827

//MAC_894 replaced by MAC_5826

//MAC_905 replaced by MAC_5827

//MAC_904 replaced by MAC_5827

//MAC_903 replaced by MAC_5826

//MAC_902 replaced by MAC_5827

//MAC_901 replaced by MAC_5827

//MAC_900 replaced by MAC_5826

//MAC_911 replaced by MAC_5827

//MAC_910 replaced by MAC_5827

//MAC_909 replaced by MAC_5826

//MAC_908 replaced by MAC_5827

//MAC_907 replaced by MAC_5827

//MAC_906 replaced by MAC_5826

//MAC_917 replaced by MAC_5827

//MAC_916 replaced by MAC_5827

//MAC_915 replaced by MAC_5826

//MAC_914 replaced by MAC_5827

//MAC_913 replaced by MAC_5827

//MAC_912 replaced by MAC_5826

//MAC_923 replaced by MAC_5827

//MAC_922 replaced by MAC_5827

//MAC_921 replaced by MAC_5826

//MAC_920 replaced by MAC_5827

//MAC_919 replaced by MAC_5827

//MAC_918 replaced by MAC_5826

//MAC_929 replaced by MAC_5827

//MAC_928 replaced by MAC_5827

//MAC_927 replaced by MAC_5826

//MAC_926 replaced by MAC_5827

//MAC_925 replaced by MAC_5827

//MAC_924 replaced by MAC_5826

//MAC_935 replaced by MAC_5827

//MAC_934 replaced by MAC_5827

//MAC_933 replaced by MAC_5826

//MAC_932 replaced by MAC_5827

//MAC_931 replaced by MAC_5827

//MAC_930 replaced by MAC_5826

//MAC_941 replaced by MAC_5827

//MAC_940 replaced by MAC_5827

//MAC_939 replaced by MAC_5826

//MAC_938 replaced by MAC_5827

//MAC_937 replaced by MAC_5827

//MAC_936 replaced by MAC_5826

//MAC_947 replaced by MAC_5827

//MAC_946 replaced by MAC_5827

//MAC_945 replaced by MAC_5826

//MAC_944 replaced by MAC_5827

//MAC_943 replaced by MAC_5827

//MAC_942 replaced by MAC_5826

//MAC_953 replaced by MAC_5827

//MAC_952 replaced by MAC_5827

//MAC_951 replaced by MAC_5826

//MAC_950 replaced by MAC_5827

//MAC_949 replaced by MAC_5827

//MAC_948 replaced by MAC_5826

//MAC_959 replaced by MAC_5827

//MAC_958 replaced by MAC_5827

//MAC_957 replaced by MAC_5826

//MAC_956 replaced by MAC_5827

//MAC_955 replaced by MAC_5827

//MAC_954 replaced by MAC_5826

//MAC_965 replaced by MAC_5827

//MAC_964 replaced by MAC_5827

//MAC_963 replaced by MAC_5826

//MAC_962 replaced by MAC_5827

//MAC_961 replaced by MAC_5827

//MAC_960 replaced by MAC_5826

//MAC_971 replaced by MAC_5827

//MAC_970 replaced by MAC_5827

//MAC_969 replaced by MAC_5826

//MAC_968 replaced by MAC_5827

//MAC_967 replaced by MAC_5827

//MAC_966 replaced by MAC_5826

//MAC_977 replaced by MAC_5827

//MAC_976 replaced by MAC_5827

//MAC_975 replaced by MAC_5826

//MAC_974 replaced by MAC_5827

//MAC_973 replaced by MAC_5827

//MAC_972 replaced by MAC_5826

//MAC_983 replaced by MAC_5827

//MAC_982 replaced by MAC_5827

//MAC_981 replaced by MAC_5826

//MAC_980 replaced by MAC_5827

//MAC_979 replaced by MAC_5827

//MAC_978 replaced by MAC_5826

//MAC_989 replaced by MAC_5827

//MAC_988 replaced by MAC_5827

//MAC_987 replaced by MAC_5826

//MAC_986 replaced by MAC_5827

//MAC_985 replaced by MAC_5827

//MAC_984 replaced by MAC_5826

//MAC_995 replaced by MAC_5827

//MAC_994 replaced by MAC_5827

//MAC_993 replaced by MAC_5826

//MAC_992 replaced by MAC_5827

//MAC_991 replaced by MAC_5827

//MAC_990 replaced by MAC_5826

//MAC_1001 replaced by MAC_5827

//MAC_1000 replaced by MAC_5827

//MAC_999 replaced by MAC_5826

//MAC_998 replaced by MAC_5827

//MAC_997 replaced by MAC_5827

//MAC_996 replaced by MAC_5826

//MAC_1007 replaced by MAC_5827

//MAC_1006 replaced by MAC_5827

//MAC_1005 replaced by MAC_5826

//MAC_1004 replaced by MAC_5827

//MAC_1003 replaced by MAC_5827

//MAC_1002 replaced by MAC_5826

//MAC_1013 replaced by MAC_5827

//MAC_1012 replaced by MAC_5827

//MAC_1011 replaced by MAC_5826

//MAC_1010 replaced by MAC_5827

//MAC_1009 replaced by MAC_5827

//MAC_1008 replaced by MAC_5826

//MAC_1019 replaced by MAC_5827

//MAC_1018 replaced by MAC_5827

//MAC_1017 replaced by MAC_5826

//MAC_1016 replaced by MAC_5827

//MAC_1015 replaced by MAC_5827

//MAC_1014 replaced by MAC_5826

//MAC_1025 replaced by MAC_5827

//MAC_1024 replaced by MAC_5827

//MAC_1023 replaced by MAC_5826

//MAC_1022 replaced by MAC_5827

//MAC_1021 replaced by MAC_5827

//MAC_1020 replaced by MAC_5826

//MAC_1031 replaced by MAC_5827

//MAC_1030 replaced by MAC_5827

//MAC_1029 replaced by MAC_5826

//MAC_1028 replaced by MAC_5827

//MAC_1027 replaced by MAC_5827

//MAC_1026 replaced by MAC_5826

//MAC_1037 replaced by MAC_5827

//MAC_1036 replaced by MAC_5827

//MAC_1035 replaced by MAC_5826

//MAC_1034 replaced by MAC_5827

//MAC_1033 replaced by MAC_5827

//MAC_1032 replaced by MAC_5826

//MAC_1043 replaced by MAC_5827

//MAC_1042 replaced by MAC_5827

//MAC_1041 replaced by MAC_5826

//MAC_1040 replaced by MAC_5827

//MAC_1039 replaced by MAC_5827

//MAC_1038 replaced by MAC_5826

//MAC_1049 replaced by MAC_5827

//MAC_1048 replaced by MAC_5827

//MAC_1047 replaced by MAC_5826

//MAC_1046 replaced by MAC_5827

//MAC_1045 replaced by MAC_5827

//MAC_1044 replaced by MAC_5826

//MAC_1055 replaced by MAC_5827

//MAC_1054 replaced by MAC_5827

//MAC_1053 replaced by MAC_5826

//MAC_1052 replaced by MAC_5827

//MAC_1051 replaced by MAC_5827

//MAC_1050 replaced by MAC_5826

//MAC_1061 replaced by MAC_5827

//MAC_1060 replaced by MAC_5827

//MAC_1059 replaced by MAC_5826

//MAC_1058 replaced by MAC_5827

//MAC_1057 replaced by MAC_5827

//MAC_1056 replaced by MAC_5826

//MAC_1067 replaced by MAC_5827

//MAC_1066 replaced by MAC_5827

//MAC_1065 replaced by MAC_5826

//MAC_1064 replaced by MAC_5827

//MAC_1063 replaced by MAC_5827

//MAC_1062 replaced by MAC_5826

//MAC_1073 replaced by MAC_5827

//MAC_1072 replaced by MAC_5827

//MAC_1071 replaced by MAC_5826

//MAC_1070 replaced by MAC_5827

//MAC_1069 replaced by MAC_5827

//MAC_1068 replaced by MAC_5826

//MAC_1079 replaced by MAC_5827

//MAC_1078 replaced by MAC_5827

//MAC_1077 replaced by MAC_5826

//MAC_1076 replaced by MAC_5827

//MAC_1075 replaced by MAC_5827

//MAC_1074 replaced by MAC_5826

//MAC_1085 replaced by MAC_5827

//MAC_1084 replaced by MAC_5827

//MAC_1083 replaced by MAC_5826

//MAC_1082 replaced by MAC_5827

//MAC_1081 replaced by MAC_5827

//MAC_1080 replaced by MAC_5826

//MAC_1091 replaced by MAC_5827

//MAC_1090 replaced by MAC_5827

//MAC_1089 replaced by MAC_5826

//MAC_1088 replaced by MAC_5827

//MAC_1087 replaced by MAC_5827

//MAC_1086 replaced by MAC_5826

//MAC_1097 replaced by MAC_5827

//MAC_1096 replaced by MAC_5827

//MAC_1095 replaced by MAC_5826

//MAC_1094 replaced by MAC_5827

//MAC_1093 replaced by MAC_5827

//MAC_1092 replaced by MAC_5826

//MAC_1103 replaced by MAC_5827

//MAC_1102 replaced by MAC_5827

//MAC_1101 replaced by MAC_5826

//MAC_1100 replaced by MAC_5827

//MAC_1099 replaced by MAC_5827

//MAC_1098 replaced by MAC_5826

//MAC_1109 replaced by MAC_5827

//MAC_1108 replaced by MAC_5827

//MAC_1107 replaced by MAC_5826

//MAC_1106 replaced by MAC_5827

//MAC_1105 replaced by MAC_5827

//MAC_1104 replaced by MAC_5826

//MAC_1115 replaced by MAC_5827

//MAC_1114 replaced by MAC_5827

//MAC_1113 replaced by MAC_5826

//MAC_1112 replaced by MAC_5827

//MAC_1111 replaced by MAC_5827

//MAC_1110 replaced by MAC_5826

//MAC_1121 replaced by MAC_5827

//MAC_1120 replaced by MAC_5827

//MAC_1119 replaced by MAC_5826

//MAC_1118 replaced by MAC_5827

//MAC_1117 replaced by MAC_5827

//MAC_1116 replaced by MAC_5826

//MAC_1127 replaced by MAC_5827

//MAC_1126 replaced by MAC_5827

//MAC_1125 replaced by MAC_5826

//MAC_1124 replaced by MAC_5827

//MAC_1123 replaced by MAC_5827

//MAC_1122 replaced by MAC_5826

//MAC_1133 replaced by MAC_5827

//MAC_1132 replaced by MAC_5827

//MAC_1131 replaced by MAC_5826

//MAC_1130 replaced by MAC_5827

//MAC_1129 replaced by MAC_5827

//MAC_1128 replaced by MAC_5826

//MAC_1139 replaced by MAC_5827

//MAC_1138 replaced by MAC_5827

//MAC_1137 replaced by MAC_5826

//MAC_1136 replaced by MAC_5827

//MAC_1135 replaced by MAC_5827

//MAC_1134 replaced by MAC_5826

//MAC_1145 replaced by MAC_5827

//MAC_1144 replaced by MAC_5827

//MAC_1143 replaced by MAC_5826

//MAC_1142 replaced by MAC_5827

//MAC_1141 replaced by MAC_5827

//MAC_1140 replaced by MAC_5826

//MAC_1151 replaced by MAC_5827

//MAC_1150 replaced by MAC_5827

//MAC_1149 replaced by MAC_5826

//MAC_1148 replaced by MAC_5827

//MAC_1147 replaced by MAC_5827

//MAC_1146 replaced by MAC_5826

//MAC_1157 replaced by MAC_5827

//MAC_1156 replaced by MAC_5827

//MAC_1155 replaced by MAC_5826

//MAC_1154 replaced by MAC_5827

//MAC_1153 replaced by MAC_5827

//MAC_1152 replaced by MAC_5826

//MAC_1163 replaced by MAC_5827

//MAC_1162 replaced by MAC_5827

//MAC_1161 replaced by MAC_5826

//MAC_1160 replaced by MAC_5827

//MAC_1159 replaced by MAC_5827

//MAC_1158 replaced by MAC_5826

//MAC_1169 replaced by MAC_5827

//MAC_1168 replaced by MAC_5827

//MAC_1167 replaced by MAC_5826

//MAC_1166 replaced by MAC_5827

//MAC_1165 replaced by MAC_5827

//MAC_1164 replaced by MAC_5826

//MAC_1175 replaced by MAC_5827

//MAC_1174 replaced by MAC_5827

//MAC_1173 replaced by MAC_5826

//MAC_1172 replaced by MAC_5827

//MAC_1171 replaced by MAC_5827

//MAC_1170 replaced by MAC_5826

//MAC_1181 replaced by MAC_5827

//MAC_1180 replaced by MAC_5827

//MAC_1179 replaced by MAC_5826

//MAC_1178 replaced by MAC_5827

//MAC_1177 replaced by MAC_5827

//MAC_1176 replaced by MAC_5826

//MAC_1187 replaced by MAC_5827

//MAC_1186 replaced by MAC_5827

//MAC_1185 replaced by MAC_5826

//MAC_1184 replaced by MAC_5827

//MAC_1183 replaced by MAC_5827

//MAC_1182 replaced by MAC_5826

//MAC_1193 replaced by MAC_5827

//MAC_1192 replaced by MAC_5827

//MAC_1191 replaced by MAC_5826

//MAC_1190 replaced by MAC_5827

//MAC_1189 replaced by MAC_5827

//MAC_1188 replaced by MAC_5826

//MAC_1199 replaced by MAC_5827

//MAC_1198 replaced by MAC_5827

//MAC_1197 replaced by MAC_5826

//MAC_1196 replaced by MAC_5827

//MAC_1195 replaced by MAC_5827

//MAC_1194 replaced by MAC_5826

//MAC_1205 replaced by MAC_5827

//MAC_1204 replaced by MAC_5827

//MAC_1203 replaced by MAC_5826

//MAC_1202 replaced by MAC_5827

//MAC_1201 replaced by MAC_5827

//MAC_1200 replaced by MAC_5826

//MAC_1211 replaced by MAC_5827

//MAC_1210 replaced by MAC_5827

//MAC_1209 replaced by MAC_5826

//MAC_1208 replaced by MAC_5827

//MAC_1207 replaced by MAC_5827

//MAC_1206 replaced by MAC_5826

//MAC_1217 replaced by MAC_5827

//MAC_1216 replaced by MAC_5827

//MAC_1215 replaced by MAC_5826

//MAC_1214 replaced by MAC_5827

//MAC_1213 replaced by MAC_5827

//MAC_1212 replaced by MAC_5826

//MAC_1223 replaced by MAC_5827

//MAC_1222 replaced by MAC_5827

//MAC_1221 replaced by MAC_5826

//MAC_1220 replaced by MAC_5827

//MAC_1219 replaced by MAC_5827

//MAC_1218 replaced by MAC_5826

//MAC_1229 replaced by MAC_5827

//MAC_1228 replaced by MAC_5827

//MAC_1227 replaced by MAC_5826

//MAC_1226 replaced by MAC_5827

//MAC_1225 replaced by MAC_5827

//MAC_1224 replaced by MAC_5826

//MAC_1235 replaced by MAC_5827

//MAC_1234 replaced by MAC_5827

//MAC_1233 replaced by MAC_5826

//MAC_1232 replaced by MAC_5827

//MAC_1231 replaced by MAC_5827

//MAC_1230 replaced by MAC_5826

//MAC_1241 replaced by MAC_5827

//MAC_1240 replaced by MAC_5827

//MAC_1239 replaced by MAC_5826

//MAC_1238 replaced by MAC_5827

//MAC_1237 replaced by MAC_5827

//MAC_1236 replaced by MAC_5826

//MAC_1247 replaced by MAC_5827

//MAC_1246 replaced by MAC_5827

//MAC_1245 replaced by MAC_5826

//MAC_1244 replaced by MAC_5827

//MAC_1243 replaced by MAC_5827

//MAC_1242 replaced by MAC_5826

//MAC_1253 replaced by MAC_5827

//MAC_1252 replaced by MAC_5827

//MAC_1251 replaced by MAC_5826

//MAC_1250 replaced by MAC_5827

//MAC_1249 replaced by MAC_5827

//MAC_1248 replaced by MAC_5826

//MAC_1259 replaced by MAC_5827

//MAC_1258 replaced by MAC_5827

//MAC_1257 replaced by MAC_5826

//MAC_1256 replaced by MAC_5827

//MAC_1255 replaced by MAC_5827

//MAC_1254 replaced by MAC_5826

//MAC_1265 replaced by MAC_5827

//MAC_1264 replaced by MAC_5827

//MAC_1263 replaced by MAC_5826

//MAC_1262 replaced by MAC_5827

//MAC_1261 replaced by MAC_5827

//MAC_1260 replaced by MAC_5826

//MAC_1271 replaced by MAC_5827

//MAC_1270 replaced by MAC_5827

//MAC_1269 replaced by MAC_5826

//MAC_1268 replaced by MAC_5827

//MAC_1267 replaced by MAC_5827

//MAC_1266 replaced by MAC_5826

//MAC_1277 replaced by MAC_5827

//MAC_1276 replaced by MAC_5827

//MAC_1275 replaced by MAC_5826

//MAC_1274 replaced by MAC_5827

//MAC_1273 replaced by MAC_5827

//MAC_1272 replaced by MAC_5826

//MAC_1283 replaced by MAC_5827

//MAC_1282 replaced by MAC_5827

//MAC_1281 replaced by MAC_5826

//MAC_1280 replaced by MAC_5827

//MAC_1279 replaced by MAC_5827

//MAC_1278 replaced by MAC_5826

//MAC_1289 replaced by MAC_5827

//MAC_1288 replaced by MAC_5827

//MAC_1287 replaced by MAC_5826

//MAC_1286 replaced by MAC_5827

//MAC_1285 replaced by MAC_5827

//MAC_1284 replaced by MAC_5826

//MAC_1295 replaced by MAC_5827

//MAC_1294 replaced by MAC_5827

//MAC_1293 replaced by MAC_5826

//MAC_1292 replaced by MAC_5827

//MAC_1291 replaced by MAC_5827

//MAC_1290 replaced by MAC_5826

//MAC_1301 replaced by MAC_5827

//MAC_1300 replaced by MAC_5827

//MAC_1299 replaced by MAC_5826

//MAC_1298 replaced by MAC_5827

//MAC_1297 replaced by MAC_5827

//MAC_1296 replaced by MAC_5826

//MAC_1307 replaced by MAC_5827

//MAC_1306 replaced by MAC_5827

//MAC_1305 replaced by MAC_5826

//MAC_1304 replaced by MAC_5827

//MAC_1303 replaced by MAC_5827

//MAC_1302 replaced by MAC_5826

//MAC_1313 replaced by MAC_5827

//MAC_1312 replaced by MAC_5827

//MAC_1311 replaced by MAC_5826

//MAC_1310 replaced by MAC_5827

//MAC_1309 replaced by MAC_5827

//MAC_1308 replaced by MAC_5826

//MAC_1319 replaced by MAC_5827

//MAC_1318 replaced by MAC_5827

//MAC_1317 replaced by MAC_5826

//MAC_1316 replaced by MAC_5827

//MAC_1315 replaced by MAC_5827

//MAC_1314 replaced by MAC_5826

//MAC_1325 replaced by MAC_5827

//MAC_1324 replaced by MAC_5827

//MAC_1323 replaced by MAC_5826

//MAC_1322 replaced by MAC_5827

//MAC_1321 replaced by MAC_5827

//MAC_1320 replaced by MAC_5826

//MAC_1331 replaced by MAC_5827

//MAC_1330 replaced by MAC_5827

//MAC_1329 replaced by MAC_5826

//MAC_1328 replaced by MAC_5827

//MAC_1327 replaced by MAC_5827

//MAC_1326 replaced by MAC_5826

//MAC_1337 replaced by MAC_5827

//MAC_1336 replaced by MAC_5827

//MAC_1335 replaced by MAC_5826

//MAC_1334 replaced by MAC_5827

//MAC_1333 replaced by MAC_5827

//MAC_1332 replaced by MAC_5826

//MAC_1343 replaced by MAC_5827

//MAC_1342 replaced by MAC_5827

//MAC_1341 replaced by MAC_5826

//MAC_1340 replaced by MAC_5827

//MAC_1339 replaced by MAC_5827

//MAC_1338 replaced by MAC_5826

//MAC_1349 replaced by MAC_5827

//MAC_1348 replaced by MAC_5827

//MAC_1347 replaced by MAC_5826

//MAC_1346 replaced by MAC_5827

//MAC_1345 replaced by MAC_5827

//MAC_1344 replaced by MAC_5826

//MAC_1355 replaced by MAC_5827

//MAC_1354 replaced by MAC_5827

//MAC_1353 replaced by MAC_5826

//MAC_1352 replaced by MAC_5827

//MAC_1351 replaced by MAC_5827

//MAC_1350 replaced by MAC_5826

//MAC_1361 replaced by MAC_5827

//MAC_1360 replaced by MAC_5827

//MAC_1359 replaced by MAC_5826

//MAC_1358 replaced by MAC_5827

//MAC_1357 replaced by MAC_5827

//MAC_1356 replaced by MAC_5826

//MAC_1367 replaced by MAC_5827

//MAC_1366 replaced by MAC_5827

//MAC_1365 replaced by MAC_5826

//MAC_1364 replaced by MAC_5827

//MAC_1363 replaced by MAC_5827

//MAC_1362 replaced by MAC_5826

//MAC_1373 replaced by MAC_5827

//MAC_1372 replaced by MAC_5827

//MAC_1371 replaced by MAC_5826

//MAC_1370 replaced by MAC_5827

//MAC_1369 replaced by MAC_5827

//MAC_1368 replaced by MAC_5826

//MAC_1379 replaced by MAC_5827

//MAC_1378 replaced by MAC_5827

//MAC_1377 replaced by MAC_5826

//MAC_1376 replaced by MAC_5827

//MAC_1375 replaced by MAC_5827

//MAC_1374 replaced by MAC_5826

//MAC_1385 replaced by MAC_5827

//MAC_1384 replaced by MAC_5827

//MAC_1383 replaced by MAC_5826

//MAC_1382 replaced by MAC_5827

//MAC_1381 replaced by MAC_5827

//MAC_1380 replaced by MAC_5826

//MAC_1391 replaced by MAC_5827

//MAC_1390 replaced by MAC_5827

//MAC_1389 replaced by MAC_5826

//MAC_1388 replaced by MAC_5827

//MAC_1387 replaced by MAC_5827

//MAC_1386 replaced by MAC_5826

//MAC_1397 replaced by MAC_5827

//MAC_1396 replaced by MAC_5827

//MAC_1395 replaced by MAC_5826

//MAC_1394 replaced by MAC_5827

//MAC_1393 replaced by MAC_5827

//MAC_1392 replaced by MAC_5826

//MAC_1403 replaced by MAC_5827

//MAC_1402 replaced by MAC_5827

//MAC_1401 replaced by MAC_5826

//MAC_1400 replaced by MAC_5827

//MAC_1399 replaced by MAC_5827

//MAC_1398 replaced by MAC_5826

//MAC_1409 replaced by MAC_5827

//MAC_1408 replaced by MAC_5827

//MAC_1407 replaced by MAC_5826

//MAC_1406 replaced by MAC_5827

//MAC_1405 replaced by MAC_5827

//MAC_1404 replaced by MAC_5826

//MAC_1415 replaced by MAC_5827

//MAC_1414 replaced by MAC_5827

//MAC_1413 replaced by MAC_5826

//MAC_1412 replaced by MAC_5827

//MAC_1411 replaced by MAC_5827

//MAC_1410 replaced by MAC_5826

//MAC_1421 replaced by MAC_5827

//MAC_1420 replaced by MAC_5827

//MAC_1419 replaced by MAC_5826

//MAC_1418 replaced by MAC_5827

//MAC_1417 replaced by MAC_5827

//MAC_1416 replaced by MAC_5826

//MAC_1427 replaced by MAC_5827

//MAC_1426 replaced by MAC_5827

//MAC_1425 replaced by MAC_5826

//MAC_1424 replaced by MAC_5827

//MAC_1423 replaced by MAC_5827

//MAC_1422 replaced by MAC_5826

//MAC_1433 replaced by MAC_5827

//MAC_1432 replaced by MAC_5827

//MAC_1431 replaced by MAC_5826

//MAC_1430 replaced by MAC_5827

//MAC_1429 replaced by MAC_5827

//MAC_1428 replaced by MAC_5826

//MAC_1439 replaced by MAC_5827

//MAC_1438 replaced by MAC_5827

//MAC_1437 replaced by MAC_5826

//MAC_1436 replaced by MAC_5827

//MAC_1435 replaced by MAC_5827

//MAC_1434 replaced by MAC_5826

//MAC_1445 replaced by MAC_5827

//MAC_1444 replaced by MAC_5827

//MAC_1443 replaced by MAC_5826

//MAC_1442 replaced by MAC_5827

//MAC_1441 replaced by MAC_5827

//MAC_1440 replaced by MAC_5826

//MAC_1451 replaced by MAC_5827

//MAC_1450 replaced by MAC_5827

//MAC_1449 replaced by MAC_5826

//MAC_1448 replaced by MAC_5827

//MAC_1447 replaced by MAC_5827

//MAC_1446 replaced by MAC_5826

//MAC_1457 replaced by MAC_5827

//MAC_1456 replaced by MAC_5827

//MAC_1455 replaced by MAC_5826

//MAC_1454 replaced by MAC_5827

//MAC_1453 replaced by MAC_5827

//MAC_1452 replaced by MAC_5826

//MAC_1463 replaced by MAC_5827

//MAC_1462 replaced by MAC_5827

//MAC_1461 replaced by MAC_5826

//MAC_1460 replaced by MAC_5827

//MAC_1459 replaced by MAC_5827

//MAC_1458 replaced by MAC_5826

//MAC_1469 replaced by MAC_5827

//MAC_1468 replaced by MAC_5827

//MAC_1467 replaced by MAC_5826

//MAC_1466 replaced by MAC_5827

//MAC_1465 replaced by MAC_5827

//MAC_1464 replaced by MAC_5826

//MAC_1475 replaced by MAC_5827

//MAC_1474 replaced by MAC_5827

//MAC_1473 replaced by MAC_5826

//MAC_1472 replaced by MAC_5827

//MAC_1471 replaced by MAC_5827

//MAC_1470 replaced by MAC_5826

//MAC_1481 replaced by MAC_5827

//MAC_1480 replaced by MAC_5827

//MAC_1479 replaced by MAC_5826

//MAC_1478 replaced by MAC_5827

//MAC_1477 replaced by MAC_5827

//MAC_1476 replaced by MAC_5826

//MAC_1487 replaced by MAC_5827

//MAC_1486 replaced by MAC_5827

//MAC_1485 replaced by MAC_5826

//MAC_1484 replaced by MAC_5827

//MAC_1483 replaced by MAC_5827

//MAC_1482 replaced by MAC_5826

//MAC_1493 replaced by MAC_5827

//MAC_1492 replaced by MAC_5827

//MAC_1491 replaced by MAC_5826

//MAC_1490 replaced by MAC_5827

//MAC_1489 replaced by MAC_5827

//MAC_1488 replaced by MAC_5826

//MAC_1499 replaced by MAC_5827

//MAC_1498 replaced by MAC_5827

//MAC_1497 replaced by MAC_5826

//MAC_1496 replaced by MAC_5827

//MAC_1495 replaced by MAC_5827

//MAC_1494 replaced by MAC_5826

//MAC_1505 replaced by MAC_5827

//MAC_1504 replaced by MAC_5827

//MAC_1503 replaced by MAC_5826

//MAC_1502 replaced by MAC_5827

//MAC_1501 replaced by MAC_5827

//MAC_1500 replaced by MAC_5826

//MAC_1511 replaced by MAC_5827

//MAC_1510 replaced by MAC_5827

//MAC_1509 replaced by MAC_5826

//MAC_1508 replaced by MAC_5827

//MAC_1507 replaced by MAC_5827

//MAC_1506 replaced by MAC_5826

//MAC_1517 replaced by MAC_5827

//MAC_1516 replaced by MAC_5827

//MAC_1515 replaced by MAC_5826

//MAC_1514 replaced by MAC_5827

//MAC_1513 replaced by MAC_5827

//MAC_1512 replaced by MAC_5826

//MAC_1523 replaced by MAC_5827

//MAC_1522 replaced by MAC_5827

//MAC_1521 replaced by MAC_5826

//MAC_1520 replaced by MAC_5827

//MAC_1519 replaced by MAC_5827

//MAC_1518 replaced by MAC_5826

//MAC_1529 replaced by MAC_5827

//MAC_1528 replaced by MAC_5827

//MAC_1527 replaced by MAC_5826

//MAC_1526 replaced by MAC_5827

//MAC_1525 replaced by MAC_5827

//MAC_1524 replaced by MAC_5826

//MAC_1535 replaced by MAC_5827

//MAC_1534 replaced by MAC_5827

//MAC_1533 replaced by MAC_5826

//MAC_1532 replaced by MAC_5827

//MAC_1531 replaced by MAC_5827

//MAC_1530 replaced by MAC_5826

//MAC_1541 replaced by MAC_5827

//MAC_1540 replaced by MAC_5827

//MAC_1539 replaced by MAC_5826

//MAC_1538 replaced by MAC_5827

//MAC_1537 replaced by MAC_5827

//MAC_1536 replaced by MAC_5826

//MAC_1547 replaced by MAC_5827

//MAC_1546 replaced by MAC_5827

//MAC_1545 replaced by MAC_5826

//MAC_1544 replaced by MAC_5827

//MAC_1543 replaced by MAC_5827

//MAC_1542 replaced by MAC_5826

//MAC_1553 replaced by MAC_5827

//MAC_1552 replaced by MAC_5827

//MAC_1551 replaced by MAC_5826

//MAC_1550 replaced by MAC_5827

//MAC_1549 replaced by MAC_5827

//MAC_1548 replaced by MAC_5826

//MAC_1559 replaced by MAC_5827

//MAC_1558 replaced by MAC_5827

//MAC_1557 replaced by MAC_5826

//MAC_1556 replaced by MAC_5827

//MAC_1555 replaced by MAC_5827

//MAC_1554 replaced by MAC_5826

//MAC_1565 replaced by MAC_5827

//MAC_1564 replaced by MAC_5827

//MAC_1563 replaced by MAC_5826

//MAC_1562 replaced by MAC_5827

//MAC_1561 replaced by MAC_5827

//MAC_1560 replaced by MAC_5826

//MAC_1571 replaced by MAC_5827

//MAC_1570 replaced by MAC_5827

//MAC_1569 replaced by MAC_5826

//MAC_1568 replaced by MAC_5827

//MAC_1567 replaced by MAC_5827

//MAC_1566 replaced by MAC_5826

//MAC_1577 replaced by MAC_5827

//MAC_1576 replaced by MAC_5827

//MAC_1575 replaced by MAC_5826

//MAC_1574 replaced by MAC_5827

//MAC_1573 replaced by MAC_5827

//MAC_1572 replaced by MAC_5826

//MAC_1583 replaced by MAC_5827

//MAC_1582 replaced by MAC_5827

//MAC_1581 replaced by MAC_5826

//MAC_1580 replaced by MAC_5827

//MAC_1579 replaced by MAC_5827

//MAC_1578 replaced by MAC_5826

//MAC_1589 replaced by MAC_5827

//MAC_1588 replaced by MAC_5827

//MAC_1587 replaced by MAC_5826

//MAC_1586 replaced by MAC_5827

//MAC_1585 replaced by MAC_5827

//MAC_1584 replaced by MAC_5826

//MAC_1595 replaced by MAC_5827

//MAC_1594 replaced by MAC_5827

//MAC_1593 replaced by MAC_5826

//MAC_1592 replaced by MAC_5827

//MAC_1591 replaced by MAC_5827

//MAC_1590 replaced by MAC_5826

//MAC_1601 replaced by MAC_5827

//MAC_1600 replaced by MAC_5827

//MAC_1599 replaced by MAC_5826

//MAC_1598 replaced by MAC_5827

//MAC_1597 replaced by MAC_5827

//MAC_1596 replaced by MAC_5826

//MAC_1607 replaced by MAC_5827

//MAC_1606 replaced by MAC_5827

//MAC_1605 replaced by MAC_5826

//MAC_1604 replaced by MAC_5827

//MAC_1603 replaced by MAC_5827

//MAC_1602 replaced by MAC_5826

//MAC_1613 replaced by MAC_5827

//MAC_1612 replaced by MAC_5827

//MAC_1611 replaced by MAC_5826

//MAC_1610 replaced by MAC_5827

//MAC_1609 replaced by MAC_5827

//MAC_1608 replaced by MAC_5826

//MAC_1619 replaced by MAC_5827

//MAC_1618 replaced by MAC_5827

//MAC_1617 replaced by MAC_5826

//MAC_1616 replaced by MAC_5827

//MAC_1615 replaced by MAC_5827

//MAC_1614 replaced by MAC_5826

//MAC_1625 replaced by MAC_5827

//MAC_1624 replaced by MAC_5827

//MAC_1623 replaced by MAC_5826

//MAC_1622 replaced by MAC_5827

//MAC_1621 replaced by MAC_5827

//MAC_1620 replaced by MAC_5826

//MAC_1631 replaced by MAC_5827

//MAC_1630 replaced by MAC_5827

//MAC_1629 replaced by MAC_5826

//MAC_1628 replaced by MAC_5827

//MAC_1627 replaced by MAC_5827

//MAC_1626 replaced by MAC_5826

//MAC_1637 replaced by MAC_5827

//MAC_1636 replaced by MAC_5827

//MAC_1635 replaced by MAC_5826

//MAC_1634 replaced by MAC_5827

//MAC_1633 replaced by MAC_5827

//MAC_1632 replaced by MAC_5826

//MAC_1643 replaced by MAC_5827

//MAC_1642 replaced by MAC_5827

//MAC_1641 replaced by MAC_5826

//MAC_1640 replaced by MAC_5827

//MAC_1639 replaced by MAC_5827

//MAC_1638 replaced by MAC_5826

//MAC_1649 replaced by MAC_5827

//MAC_1648 replaced by MAC_5827

//MAC_1647 replaced by MAC_5826

//MAC_1646 replaced by MAC_5827

//MAC_1645 replaced by MAC_5827

//MAC_1644 replaced by MAC_5826

//MAC_1655 replaced by MAC_5827

//MAC_1654 replaced by MAC_5827

//MAC_1653 replaced by MAC_5826

//MAC_1652 replaced by MAC_5827

//MAC_1651 replaced by MAC_5827

//MAC_1650 replaced by MAC_5826

//MAC_1661 replaced by MAC_5827

//MAC_1660 replaced by MAC_5827

//MAC_1659 replaced by MAC_5826

//MAC_1658 replaced by MAC_5827

//MAC_1657 replaced by MAC_5827

//MAC_1656 replaced by MAC_5826

//MAC_1667 replaced by MAC_5827

//MAC_1666 replaced by MAC_5827

//MAC_1665 replaced by MAC_5826

//MAC_1664 replaced by MAC_5827

//MAC_1663 replaced by MAC_5827

//MAC_1662 replaced by MAC_5826

//MAC_1673 replaced by MAC_5827

//MAC_1672 replaced by MAC_5827

//MAC_1671 replaced by MAC_5826

//MAC_1670 replaced by MAC_5827

//MAC_1669 replaced by MAC_5827

//MAC_1668 replaced by MAC_5826

//MAC_1679 replaced by MAC_5827

//MAC_1678 replaced by MAC_5827

//MAC_1677 replaced by MAC_5826

//MAC_1676 replaced by MAC_5827

//MAC_1675 replaced by MAC_5827

//MAC_1674 replaced by MAC_5826

//MAC_1685 replaced by MAC_5827

//MAC_1684 replaced by MAC_5827

//MAC_1683 replaced by MAC_5826

//MAC_1682 replaced by MAC_5827

//MAC_1681 replaced by MAC_5827

//MAC_1680 replaced by MAC_5826

//MAC_1691 replaced by MAC_5827

//MAC_1690 replaced by MAC_5827

//MAC_1689 replaced by MAC_5826

//MAC_1688 replaced by MAC_5827

//MAC_1687 replaced by MAC_5827

//MAC_1686 replaced by MAC_5826

//MAC_1697 replaced by MAC_5827

//MAC_1696 replaced by MAC_5827

//MAC_1695 replaced by MAC_5826

//MAC_1694 replaced by MAC_5827

//MAC_1693 replaced by MAC_5827

//MAC_1692 replaced by MAC_5826

//MAC_1703 replaced by MAC_5827

//MAC_1702 replaced by MAC_5827

//MAC_1701 replaced by MAC_5826

//MAC_1700 replaced by MAC_5827

//MAC_1699 replaced by MAC_5827

//MAC_1698 replaced by MAC_5826

//MAC_1709 replaced by MAC_5827

//MAC_1708 replaced by MAC_5827

//MAC_1707 replaced by MAC_5826

//MAC_1706 replaced by MAC_5827

//MAC_1705 replaced by MAC_5827

//MAC_1704 replaced by MAC_5826

//MAC_1715 replaced by MAC_5827

//MAC_1714 replaced by MAC_5827

//MAC_1713 replaced by MAC_5826

//MAC_1712 replaced by MAC_5827

//MAC_1711 replaced by MAC_5827

//MAC_1710 replaced by MAC_5826

//MAC_1721 replaced by MAC_5827

//MAC_1720 replaced by MAC_5827

//MAC_1719 replaced by MAC_5826

//MAC_1718 replaced by MAC_5827

//MAC_1717 replaced by MAC_5827

//MAC_1716 replaced by MAC_5826

//MAC_1727 replaced by MAC_5827

//MAC_1726 replaced by MAC_5827

//MAC_1725 replaced by MAC_5826

//MAC_1724 replaced by MAC_5827

//MAC_1723 replaced by MAC_5827

//MAC_1722 replaced by MAC_5826

//MAC_1733 replaced by MAC_5827

//MAC_1732 replaced by MAC_5827

//MAC_1731 replaced by MAC_5826

//MAC_1730 replaced by MAC_5827

//MAC_1729 replaced by MAC_5827

//MAC_1728 replaced by MAC_5826

//MAC_1739 replaced by MAC_5827

//MAC_1738 replaced by MAC_5827

//MAC_1737 replaced by MAC_5826

//MAC_1736 replaced by MAC_5827

//MAC_1735 replaced by MAC_5827

//MAC_1734 replaced by MAC_5826

//MAC_1745 replaced by MAC_5827

//MAC_1744 replaced by MAC_5827

//MAC_1743 replaced by MAC_5826

//MAC_1742 replaced by MAC_5827

//MAC_1741 replaced by MAC_5827

//MAC_1740 replaced by MAC_5826

//MAC_1751 replaced by MAC_5827

//MAC_1750 replaced by MAC_5827

//MAC_1749 replaced by MAC_5826

//MAC_1748 replaced by MAC_5827

//MAC_1747 replaced by MAC_5827

//MAC_1746 replaced by MAC_5826

//MAC_1757 replaced by MAC_5827

//MAC_1756 replaced by MAC_5827

//MAC_1755 replaced by MAC_5826

//MAC_1754 replaced by MAC_5827

//MAC_1753 replaced by MAC_5827

//MAC_1752 replaced by MAC_5826

//MAC_1763 replaced by MAC_5827

//MAC_1762 replaced by MAC_5827

//MAC_1761 replaced by MAC_5826

//MAC_1760 replaced by MAC_5827

//MAC_1759 replaced by MAC_5827

//MAC_1758 replaced by MAC_5826

//MAC_1769 replaced by MAC_5827

//MAC_1768 replaced by MAC_5827

//MAC_1767 replaced by MAC_5826

//MAC_1766 replaced by MAC_5827

//MAC_1765 replaced by MAC_5827

//MAC_1764 replaced by MAC_5826

//MAC_1775 replaced by MAC_5827

//MAC_1774 replaced by MAC_5827

//MAC_1773 replaced by MAC_5826

//MAC_1772 replaced by MAC_5827

//MAC_1771 replaced by MAC_5827

//MAC_1770 replaced by MAC_5826

//MAC_1781 replaced by MAC_5827

//MAC_1780 replaced by MAC_5827

//MAC_1779 replaced by MAC_5826

//MAC_1778 replaced by MAC_5827

//MAC_1777 replaced by MAC_5827

//MAC_1776 replaced by MAC_5826

//MAC_1787 replaced by MAC_5827

//MAC_1786 replaced by MAC_5827

//MAC_1785 replaced by MAC_5826

//MAC_1784 replaced by MAC_5827

//MAC_1783 replaced by MAC_5827

//MAC_1782 replaced by MAC_5826

//MAC_1793 replaced by MAC_5827

//MAC_1792 replaced by MAC_5827

//MAC_1791 replaced by MAC_5826

//MAC_1790 replaced by MAC_5827

//MAC_1789 replaced by MAC_5827

//MAC_1788 replaced by MAC_5826

//MAC_1799 replaced by MAC_5827

//MAC_1798 replaced by MAC_5827

//MAC_1797 replaced by MAC_5826

//MAC_1796 replaced by MAC_5827

//MAC_1795 replaced by MAC_5827

//MAC_1794 replaced by MAC_5826

//MAC_1805 replaced by MAC_5827

//MAC_1804 replaced by MAC_5827

//MAC_1803 replaced by MAC_5826

//MAC_1802 replaced by MAC_5827

//MAC_1801 replaced by MAC_5827

//MAC_1800 replaced by MAC_5826

//MAC_1811 replaced by MAC_5827

//MAC_1810 replaced by MAC_5827

//MAC_1809 replaced by MAC_5826

//MAC_1808 replaced by MAC_5827

//MAC_1807 replaced by MAC_5827

//MAC_1806 replaced by MAC_5826

//MAC_1817 replaced by MAC_5827

//MAC_1816 replaced by MAC_5827

//MAC_1815 replaced by MAC_5826

//MAC_1814 replaced by MAC_5827

//MAC_1813 replaced by MAC_5827

//MAC_1812 replaced by MAC_5826

//MAC_1823 replaced by MAC_5827

//MAC_1822 replaced by MAC_5827

//MAC_1821 replaced by MAC_5826

//MAC_1820 replaced by MAC_5827

//MAC_1819 replaced by MAC_5827

//MAC_1818 replaced by MAC_5826

//MAC_1829 replaced by MAC_5827

//MAC_1828 replaced by MAC_5827

//MAC_1827 replaced by MAC_5826

//MAC_1826 replaced by MAC_5827

//MAC_1825 replaced by MAC_5827

//MAC_1824 replaced by MAC_5826

//MAC_1835 replaced by MAC_5827

//MAC_1834 replaced by MAC_5827

//MAC_1833 replaced by MAC_5826

//MAC_1832 replaced by MAC_5827

//MAC_1831 replaced by MAC_5827

//MAC_1830 replaced by MAC_5826

//MAC_1841 replaced by MAC_5827

//MAC_1840 replaced by MAC_5827

//MAC_1839 replaced by MAC_5826

//MAC_1838 replaced by MAC_5827

//MAC_1837 replaced by MAC_5827

//MAC_1836 replaced by MAC_5826

//MAC_1847 replaced by MAC_5827

//MAC_1846 replaced by MAC_5827

//MAC_1845 replaced by MAC_5826

//MAC_1844 replaced by MAC_5827

//MAC_1843 replaced by MAC_5827

//MAC_1842 replaced by MAC_5826

//MAC_1853 replaced by MAC_5827

//MAC_1852 replaced by MAC_5827

//MAC_1851 replaced by MAC_5826

//MAC_1850 replaced by MAC_5827

//MAC_1849 replaced by MAC_5827

//MAC_1848 replaced by MAC_5826

//MAC_1859 replaced by MAC_5827

//MAC_1858 replaced by MAC_5827

//MAC_1857 replaced by MAC_5826

//MAC_1856 replaced by MAC_5827

//MAC_1855 replaced by MAC_5827

//MAC_1854 replaced by MAC_5826

//MAC_1865 replaced by MAC_5827

//MAC_1864 replaced by MAC_5827

//MAC_1863 replaced by MAC_5826

//MAC_1862 replaced by MAC_5827

//MAC_1861 replaced by MAC_5827

//MAC_1860 replaced by MAC_5826

//MAC_1871 replaced by MAC_5827

//MAC_1870 replaced by MAC_5827

//MAC_1869 replaced by MAC_5826

//MAC_1868 replaced by MAC_5827

//MAC_1867 replaced by MAC_5827

//MAC_1866 replaced by MAC_5826

//MAC_1877 replaced by MAC_5827

//MAC_1876 replaced by MAC_5827

//MAC_1875 replaced by MAC_5826

//MAC_1874 replaced by MAC_5827

//MAC_1873 replaced by MAC_5827

//MAC_1872 replaced by MAC_5826

//MAC_1883 replaced by MAC_5827

//MAC_1882 replaced by MAC_5827

//MAC_1881 replaced by MAC_5826

//MAC_1880 replaced by MAC_5827

//MAC_1879 replaced by MAC_5827

//MAC_1878 replaced by MAC_5826

//MAC_1889 replaced by MAC_5827

//MAC_1888 replaced by MAC_5827

//MAC_1887 replaced by MAC_5826

//MAC_1886 replaced by MAC_5827

//MAC_1885 replaced by MAC_5827

//MAC_1884 replaced by MAC_5826

//MAC_1895 replaced by MAC_5827

//MAC_1894 replaced by MAC_5827

//MAC_1893 replaced by MAC_5826

//MAC_1892 replaced by MAC_5827

//MAC_1891 replaced by MAC_5827

//MAC_1890 replaced by MAC_5826

//MAC_1901 replaced by MAC_5827

//MAC_1900 replaced by MAC_5827

//MAC_1899 replaced by MAC_5826

//MAC_1898 replaced by MAC_5827

//MAC_1897 replaced by MAC_5827

//MAC_1896 replaced by MAC_5826

//MAC_1907 replaced by MAC_5827

//MAC_1906 replaced by MAC_5827

//MAC_1905 replaced by MAC_5826

//MAC_1904 replaced by MAC_5827

//MAC_1903 replaced by MAC_5827

//MAC_1902 replaced by MAC_5826

//MAC_1913 replaced by MAC_5827

//MAC_1912 replaced by MAC_5827

//MAC_1911 replaced by MAC_5826

//MAC_1910 replaced by MAC_5827

//MAC_1909 replaced by MAC_5827

//MAC_1908 replaced by MAC_5826

//MAC_1919 replaced by MAC_5827

//MAC_1918 replaced by MAC_5827

//MAC_1917 replaced by MAC_5826

//MAC_1916 replaced by MAC_5827

//MAC_1915 replaced by MAC_5827

//MAC_1914 replaced by MAC_5826

//MAC_1925 replaced by MAC_5827

//MAC_1924 replaced by MAC_5827

//MAC_1923 replaced by MAC_5826

//MAC_1922 replaced by MAC_5827

//MAC_1921 replaced by MAC_5827

//MAC_1920 replaced by MAC_5826

//MAC_1931 replaced by MAC_5827

//MAC_1930 replaced by MAC_5827

//MAC_1929 replaced by MAC_5826

//MAC_1928 replaced by MAC_5827

//MAC_1927 replaced by MAC_5827

//MAC_1926 replaced by MAC_5826

//MAC_1937 replaced by MAC_5827

//MAC_1936 replaced by MAC_5827

//MAC_1935 replaced by MAC_5826

//MAC_1934 replaced by MAC_5827

//MAC_1933 replaced by MAC_5827

//MAC_1932 replaced by MAC_5826

//MAC_1943 replaced by MAC_5827

//MAC_1942 replaced by MAC_5827

//MAC_1941 replaced by MAC_5826

//MAC_1940 replaced by MAC_5827

//MAC_1939 replaced by MAC_5827

//MAC_1938 replaced by MAC_5826

//MAC_1949 replaced by MAC_5827

//MAC_1948 replaced by MAC_5827

//MAC_1947 replaced by MAC_5826

//MAC_1946 replaced by MAC_5827

//MAC_1945 replaced by MAC_5827

//MAC_1944 replaced by MAC_5826

//MAC_1955 replaced by MAC_5827

//MAC_1954 replaced by MAC_5827

//MAC_1953 replaced by MAC_5826

//MAC_1952 replaced by MAC_5827

//MAC_1951 replaced by MAC_5827

//MAC_1950 replaced by MAC_5826

//MAC_1961 replaced by MAC_5827

//MAC_1960 replaced by MAC_5827

//MAC_1959 replaced by MAC_5826

//MAC_1958 replaced by MAC_5827

//MAC_1957 replaced by MAC_5827

//MAC_1956 replaced by MAC_5826

//MAC_1967 replaced by MAC_5827

//MAC_1966 replaced by MAC_5827

//MAC_1965 replaced by MAC_5826

//MAC_1964 replaced by MAC_5827

//MAC_1963 replaced by MAC_5827

//MAC_1962 replaced by MAC_5826

//MAC_1973 replaced by MAC_5827

//MAC_1972 replaced by MAC_5827

//MAC_1971 replaced by MAC_5826

//MAC_1970 replaced by MAC_5827

//MAC_1969 replaced by MAC_5827

//MAC_1968 replaced by MAC_5826

//MAC_1979 replaced by MAC_5827

//MAC_1978 replaced by MAC_5827

//MAC_1977 replaced by MAC_5826

//MAC_1976 replaced by MAC_5827

//MAC_1975 replaced by MAC_5827

//MAC_1974 replaced by MAC_5826

//MAC_1985 replaced by MAC_5827

//MAC_1984 replaced by MAC_5827

//MAC_1983 replaced by MAC_5826

//MAC_1982 replaced by MAC_5827

//MAC_1981 replaced by MAC_5827

//MAC_1980 replaced by MAC_5826

//MAC_1991 replaced by MAC_5827

//MAC_1990 replaced by MAC_5827

//MAC_1989 replaced by MAC_5826

//MAC_1988 replaced by MAC_5827

//MAC_1987 replaced by MAC_5827

//MAC_1986 replaced by MAC_5826

//MAC_1997 replaced by MAC_5827

//MAC_1996 replaced by MAC_5827

//MAC_1995 replaced by MAC_5826

//MAC_1994 replaced by MAC_5827

//MAC_1993 replaced by MAC_5827

//MAC_1992 replaced by MAC_5826

//MAC_2003 replaced by MAC_5827

//MAC_2002 replaced by MAC_5827

//MAC_2001 replaced by MAC_5826

//MAC_2000 replaced by MAC_5827

//MAC_1999 replaced by MAC_5827

//MAC_1998 replaced by MAC_5826

//MAC_2009 replaced by MAC_5827

//MAC_2008 replaced by MAC_5827

//MAC_2007 replaced by MAC_5826

//MAC_2006 replaced by MAC_5827

//MAC_2005 replaced by MAC_5827

//MAC_2004 replaced by MAC_5826

//MAC_2015 replaced by MAC_5827

//MAC_2014 replaced by MAC_5827

//MAC_2013 replaced by MAC_5826

//MAC_2012 replaced by MAC_5827

//MAC_2011 replaced by MAC_5827

//MAC_2010 replaced by MAC_5826

//MAC_2021 replaced by MAC_5827

//MAC_2020 replaced by MAC_5827

//MAC_2019 replaced by MAC_5826

//MAC_2018 replaced by MAC_5827

//MAC_2017 replaced by MAC_5827

//MAC_2016 replaced by MAC_5826

//MAC_2027 replaced by MAC_5827

//MAC_2026 replaced by MAC_5827

//MAC_2025 replaced by MAC_5826

//MAC_2024 replaced by MAC_5827

//MAC_2023 replaced by MAC_5827

//MAC_2022 replaced by MAC_5826

//MAC_2033 replaced by MAC_5827

//MAC_2032 replaced by MAC_5827

//MAC_2031 replaced by MAC_5826

//MAC_2030 replaced by MAC_5827

//MAC_2029 replaced by MAC_5827

//MAC_2028 replaced by MAC_5826

//MAC_2039 replaced by MAC_5827

//MAC_2038 replaced by MAC_5827

//MAC_2037 replaced by MAC_5826

//MAC_2036 replaced by MAC_5827

//MAC_2035 replaced by MAC_5827

//MAC_2034 replaced by MAC_5826

//MAC_2045 replaced by MAC_5827

//MAC_2044 replaced by MAC_5827

//MAC_2043 replaced by MAC_5826

//MAC_2042 replaced by MAC_5827

//MAC_2041 replaced by MAC_5827

//MAC_2040 replaced by MAC_5826

//MAC_2051 replaced by MAC_5827

//MAC_2050 replaced by MAC_5827

//MAC_2049 replaced by MAC_5826

//MAC_2048 replaced by MAC_5827

//MAC_2047 replaced by MAC_5827

//MAC_2046 replaced by MAC_5826

//MAC_2057 replaced by MAC_5827

//MAC_2056 replaced by MAC_5827

//MAC_2055 replaced by MAC_5826

//MAC_2054 replaced by MAC_5827

//MAC_2053 replaced by MAC_5827

//MAC_2052 replaced by MAC_5826

//MAC_2063 replaced by MAC_5827

//MAC_2062 replaced by MAC_5827

//MAC_2061 replaced by MAC_5826

//MAC_2060 replaced by MAC_5827

//MAC_2059 replaced by MAC_5827

//MAC_2058 replaced by MAC_5826

//MAC_2069 replaced by MAC_5827

//MAC_2068 replaced by MAC_5827

//MAC_2067 replaced by MAC_5826

//MAC_2066 replaced by MAC_5827

//MAC_2065 replaced by MAC_5827

//MAC_2064 replaced by MAC_5826

//MAC_2075 replaced by MAC_5827

//MAC_2074 replaced by MAC_5827

//MAC_2073 replaced by MAC_5826

//MAC_2072 replaced by MAC_5827

//MAC_2071 replaced by MAC_5827

//MAC_2070 replaced by MAC_5826

//MAC_2081 replaced by MAC_5827

//MAC_2080 replaced by MAC_5827

//MAC_2079 replaced by MAC_5826

//MAC_2078 replaced by MAC_5827

//MAC_2077 replaced by MAC_5827

//MAC_2076 replaced by MAC_5826

//MAC_2087 replaced by MAC_5827

//MAC_2086 replaced by MAC_5827

//MAC_2085 replaced by MAC_5826

//MAC_2084 replaced by MAC_5827

//MAC_2083 replaced by MAC_5827

//MAC_2082 replaced by MAC_5826

//MAC_2093 replaced by MAC_5827

//MAC_2092 replaced by MAC_5827

//MAC_2091 replaced by MAC_5826

//MAC_2090 replaced by MAC_5827

//MAC_2089 replaced by MAC_5827

//MAC_2088 replaced by MAC_5826

//MAC_2099 replaced by MAC_5827

//MAC_2098 replaced by MAC_5827

//MAC_2097 replaced by MAC_5826

//MAC_2096 replaced by MAC_5827

//MAC_2095 replaced by MAC_5827

//MAC_2094 replaced by MAC_5826

//MAC_2105 replaced by MAC_5827

//MAC_2104 replaced by MAC_5827

//MAC_2103 replaced by MAC_5826

//MAC_2102 replaced by MAC_5827

//MAC_2101 replaced by MAC_5827

//MAC_2100 replaced by MAC_5826

//MAC_2111 replaced by MAC_5827

//MAC_2110 replaced by MAC_5827

//MAC_2109 replaced by MAC_5826

//MAC_2108 replaced by MAC_5827

//MAC_2107 replaced by MAC_5827

//MAC_2106 replaced by MAC_5826

//MAC_2117 replaced by MAC_5827

//MAC_2116 replaced by MAC_5827

//MAC_2115 replaced by MAC_5826

//MAC_2114 replaced by MAC_5827

//MAC_2113 replaced by MAC_5827

//MAC_2112 replaced by MAC_5826

//MAC_2123 replaced by MAC_5827

//MAC_2122 replaced by MAC_5827

//MAC_2121 replaced by MAC_5826

//MAC_2120 replaced by MAC_5827

//MAC_2119 replaced by MAC_5827

//MAC_2118 replaced by MAC_5826

//MAC_2129 replaced by MAC_5827

//MAC_2128 replaced by MAC_5827

//MAC_2127 replaced by MAC_5826

//MAC_2126 replaced by MAC_5827

//MAC_2125 replaced by MAC_5827

//MAC_2124 replaced by MAC_5826

//MAC_2135 replaced by MAC_5827

//MAC_2134 replaced by MAC_5827

//MAC_2133 replaced by MAC_5826

//MAC_2132 replaced by MAC_5827

//MAC_2131 replaced by MAC_5827

//MAC_2130 replaced by MAC_5826

//MAC_2141 replaced by MAC_5827

//MAC_2140 replaced by MAC_5827

//MAC_2139 replaced by MAC_5826

//MAC_2138 replaced by MAC_5827

//MAC_2137 replaced by MAC_5827

//MAC_2136 replaced by MAC_5826

//MAC_2147 replaced by MAC_5827

//MAC_2146 replaced by MAC_5827

//MAC_2145 replaced by MAC_5826

//MAC_2144 replaced by MAC_5827

//MAC_2143 replaced by MAC_5827

//MAC_2142 replaced by MAC_5826

//MAC_2153 replaced by MAC_5827

//MAC_2152 replaced by MAC_5827

//MAC_2151 replaced by MAC_5826

//MAC_2150 replaced by MAC_5827

//MAC_2149 replaced by MAC_5827

//MAC_2148 replaced by MAC_5826

//MAC_2159 replaced by MAC_5827

//MAC_2158 replaced by MAC_5827

//MAC_2157 replaced by MAC_5826

//MAC_2156 replaced by MAC_5827

//MAC_2155 replaced by MAC_5827

//MAC_2154 replaced by MAC_5826

//MAC_2165 replaced by MAC_5827

//MAC_2164 replaced by MAC_5827

//MAC_2163 replaced by MAC_5826

//MAC_2162 replaced by MAC_5827

//MAC_2161 replaced by MAC_5827

//MAC_2160 replaced by MAC_5826

//MAC_2171 replaced by MAC_5827

//MAC_2170 replaced by MAC_5827

//MAC_2169 replaced by MAC_5826

//MAC_2168 replaced by MAC_5827

//MAC_2167 replaced by MAC_5827

//MAC_2166 replaced by MAC_5826

//MAC_2177 replaced by MAC_5827

//MAC_2176 replaced by MAC_5827

//MAC_2175 replaced by MAC_5826

//MAC_2174 replaced by MAC_5827

//MAC_2173 replaced by MAC_5827

//MAC_2172 replaced by MAC_5826

//MAC_2183 replaced by MAC_5827

//MAC_2182 replaced by MAC_5827

//MAC_2181 replaced by MAC_5826

//MAC_2180 replaced by MAC_5827

//MAC_2179 replaced by MAC_5827

//MAC_2178 replaced by MAC_5826

//MAC_2189 replaced by MAC_5827

//MAC_2188 replaced by MAC_5827

//MAC_2187 replaced by MAC_5826

//MAC_2186 replaced by MAC_5827

//MAC_2185 replaced by MAC_5827

//MAC_2184 replaced by MAC_5826

//MAC_2195 replaced by MAC_5827

//MAC_2194 replaced by MAC_5827

//MAC_2193 replaced by MAC_5826

//MAC_2192 replaced by MAC_5827

//MAC_2191 replaced by MAC_5827

//MAC_2190 replaced by MAC_5826

//MAC_2201 replaced by MAC_5827

//MAC_2200 replaced by MAC_5827

//MAC_2199 replaced by MAC_5826

//MAC_2198 replaced by MAC_5827

//MAC_2197 replaced by MAC_5827

//MAC_2196 replaced by MAC_5826

//MAC_2207 replaced by MAC_5827

//MAC_2206 replaced by MAC_5827

//MAC_2205 replaced by MAC_5826

//MAC_2204 replaced by MAC_5827

//MAC_2203 replaced by MAC_5827

//MAC_2202 replaced by MAC_5826

//MAC_2213 replaced by MAC_5827

//MAC_2212 replaced by MAC_5827

//MAC_2211 replaced by MAC_5826

//MAC_2210 replaced by MAC_5827

//MAC_2209 replaced by MAC_5827

//MAC_2208 replaced by MAC_5826

//MAC_2219 replaced by MAC_5827

//MAC_2218 replaced by MAC_5827

//MAC_2217 replaced by MAC_5826

//MAC_2216 replaced by MAC_5827

//MAC_2215 replaced by MAC_5827

//MAC_2214 replaced by MAC_5826

//MAC_2225 replaced by MAC_5827

//MAC_2224 replaced by MAC_5827

//MAC_2223 replaced by MAC_5826

//MAC_2222 replaced by MAC_5827

//MAC_2221 replaced by MAC_5827

//MAC_2220 replaced by MAC_5826

//MAC_2231 replaced by MAC_5827

//MAC_2230 replaced by MAC_5827

//MAC_2229 replaced by MAC_5826

//MAC_2228 replaced by MAC_5827

//MAC_2227 replaced by MAC_5827

//MAC_2226 replaced by MAC_5826

//MAC_2237 replaced by MAC_5827

//MAC_2236 replaced by MAC_5827

//MAC_2235 replaced by MAC_5826

//MAC_2234 replaced by MAC_5827

//MAC_2233 replaced by MAC_5827

//MAC_2232 replaced by MAC_5826

//MAC_2243 replaced by MAC_5827

//MAC_2242 replaced by MAC_5827

//MAC_2241 replaced by MAC_5826

//MAC_2240 replaced by MAC_5827

//MAC_2239 replaced by MAC_5827

//MAC_2238 replaced by MAC_5826

//MAC_2249 replaced by MAC_5827

//MAC_2248 replaced by MAC_5827

//MAC_2247 replaced by MAC_5826

//MAC_2246 replaced by MAC_5827

//MAC_2245 replaced by MAC_5827

//MAC_2244 replaced by MAC_5826

//MAC_2255 replaced by MAC_5827

//MAC_2254 replaced by MAC_5827

//MAC_2253 replaced by MAC_5826

//MAC_2252 replaced by MAC_5827

//MAC_2251 replaced by MAC_5827

//MAC_2250 replaced by MAC_5826

//MAC_2261 replaced by MAC_5827

//MAC_2260 replaced by MAC_5827

//MAC_2259 replaced by MAC_5826

//MAC_2258 replaced by MAC_5827

//MAC_2257 replaced by MAC_5827

//MAC_2256 replaced by MAC_5826

//MAC_2267 replaced by MAC_5827

//MAC_2266 replaced by MAC_5827

//MAC_2265 replaced by MAC_5826

//MAC_2264 replaced by MAC_5827

//MAC_2263 replaced by MAC_5827

//MAC_2262 replaced by MAC_5826

//MAC_2273 replaced by MAC_5827

//MAC_2272 replaced by MAC_5827

//MAC_2271 replaced by MAC_5826

//MAC_2270 replaced by MAC_5827

//MAC_2269 replaced by MAC_5827

//MAC_2268 replaced by MAC_5826

//MAC_2279 replaced by MAC_5827

//MAC_2278 replaced by MAC_5827

//MAC_2277 replaced by MAC_5826

//MAC_2276 replaced by MAC_5827

//MAC_2275 replaced by MAC_5827

//MAC_2274 replaced by MAC_5826

//MAC_2285 replaced by MAC_5827

//MAC_2284 replaced by MAC_5827

//MAC_2283 replaced by MAC_5826

//MAC_2282 replaced by MAC_5827

//MAC_2281 replaced by MAC_5827

//MAC_2280 replaced by MAC_5826

//MAC_2291 replaced by MAC_5827

//MAC_2290 replaced by MAC_5827

//MAC_2289 replaced by MAC_5826

//MAC_2288 replaced by MAC_5827

//MAC_2287 replaced by MAC_5827

//MAC_2286 replaced by MAC_5826

//MAC_2297 replaced by MAC_5827

//MAC_2296 replaced by MAC_5827

//MAC_2295 replaced by MAC_5826

//MAC_2294 replaced by MAC_5827

//MAC_2293 replaced by MAC_5827

//MAC_2292 replaced by MAC_5826

//MAC_2303 replaced by MAC_5827

//MAC_2302 replaced by MAC_5827

//MAC_2301 replaced by MAC_5826

//MAC_2300 replaced by MAC_5827

//MAC_2299 replaced by MAC_5827

//MAC_2298 replaced by MAC_5826

//MAC_2309 replaced by MAC_5827

//MAC_2308 replaced by MAC_5827

//MAC_2307 replaced by MAC_5826

//MAC_2306 replaced by MAC_5827

//MAC_2305 replaced by MAC_5827

//MAC_2304 replaced by MAC_5826

//MAC_2315 replaced by MAC_5827

//MAC_2314 replaced by MAC_5827

//MAC_2313 replaced by MAC_5826

//MAC_2312 replaced by MAC_5827

//MAC_2311 replaced by MAC_5827

//MAC_2310 replaced by MAC_5826

//MAC_2321 replaced by MAC_5827

//MAC_2320 replaced by MAC_5827

//MAC_2319 replaced by MAC_5826

//MAC_2318 replaced by MAC_5827

//MAC_2317 replaced by MAC_5827

//MAC_2316 replaced by MAC_5826

//MAC_2327 replaced by MAC_5827

//MAC_2326 replaced by MAC_5827

//MAC_2325 replaced by MAC_5826

//MAC_2324 replaced by MAC_5827

//MAC_2323 replaced by MAC_5827

//MAC_2322 replaced by MAC_5826

//MAC_2333 replaced by MAC_5827

//MAC_2332 replaced by MAC_5827

//MAC_2331 replaced by MAC_5826

//MAC_2330 replaced by MAC_5827

//MAC_2329 replaced by MAC_5827

//MAC_2328 replaced by MAC_5826

//MAC_2339 replaced by MAC_5827

//MAC_2338 replaced by MAC_5827

//MAC_2337 replaced by MAC_5826

//MAC_2336 replaced by MAC_5827

//MAC_2335 replaced by MAC_5827

//MAC_2334 replaced by MAC_5826

//MAC_2345 replaced by MAC_5827

//MAC_2344 replaced by MAC_5827

//MAC_2343 replaced by MAC_5826

//MAC_2342 replaced by MAC_5827

//MAC_2341 replaced by MAC_5827

//MAC_2340 replaced by MAC_5826

//MAC_2351 replaced by MAC_5827

//MAC_2350 replaced by MAC_5827

//MAC_2349 replaced by MAC_5826

//MAC_2348 replaced by MAC_5827

//MAC_2347 replaced by MAC_5827

//MAC_2346 replaced by MAC_5826

//MAC_2357 replaced by MAC_5827

//MAC_2356 replaced by MAC_5827

//MAC_2355 replaced by MAC_5826

//MAC_2354 replaced by MAC_5827

//MAC_2353 replaced by MAC_5827

//MAC_2352 replaced by MAC_5826

//MAC_2363 replaced by MAC_5827

//MAC_2362 replaced by MAC_5827

//MAC_2361 replaced by MAC_5826

//MAC_2360 replaced by MAC_5827

//MAC_2359 replaced by MAC_5827

//MAC_2358 replaced by MAC_5826

//MAC_2369 replaced by MAC_5827

//MAC_2368 replaced by MAC_5827

//MAC_2367 replaced by MAC_5826

//MAC_2366 replaced by MAC_5827

//MAC_2365 replaced by MAC_5827

//MAC_2364 replaced by MAC_5826

//MAC_2375 replaced by MAC_5827

//MAC_2374 replaced by MAC_5827

//MAC_2373 replaced by MAC_5826

//MAC_2372 replaced by MAC_5827

//MAC_2371 replaced by MAC_5827

//MAC_2370 replaced by MAC_5826

//MAC_2381 replaced by MAC_5827

//MAC_2380 replaced by MAC_5827

//MAC_2379 replaced by MAC_5826

//MAC_2378 replaced by MAC_5827

//MAC_2377 replaced by MAC_5827

//MAC_2376 replaced by MAC_5826

//MAC_2387 replaced by MAC_5827

//MAC_2386 replaced by MAC_5827

//MAC_2385 replaced by MAC_5826

//MAC_2384 replaced by MAC_5827

//MAC_2383 replaced by MAC_5827

//MAC_2382 replaced by MAC_5826

//MAC_2393 replaced by MAC_5827

//MAC_2392 replaced by MAC_5827

//MAC_2391 replaced by MAC_5826

//MAC_2390 replaced by MAC_5827

//MAC_2389 replaced by MAC_5827

//MAC_2388 replaced by MAC_5826

//MAC_2399 replaced by MAC_5827

//MAC_2398 replaced by MAC_5827

//MAC_2397 replaced by MAC_5826

//MAC_2396 replaced by MAC_5827

//MAC_2395 replaced by MAC_5827

//MAC_2394 replaced by MAC_5826

//MAC_2405 replaced by MAC_5827

//MAC_2404 replaced by MAC_5827

//MAC_2403 replaced by MAC_5826

//MAC_2402 replaced by MAC_5827

//MAC_2401 replaced by MAC_5827

//MAC_2400 replaced by MAC_5826

//MAC_2411 replaced by MAC_5827

//MAC_2410 replaced by MAC_5827

//MAC_2409 replaced by MAC_5826

//MAC_2408 replaced by MAC_5827

//MAC_2407 replaced by MAC_5827

//MAC_2406 replaced by MAC_5826

//MAC_2417 replaced by MAC_5827

//MAC_2416 replaced by MAC_5827

//MAC_2415 replaced by MAC_5826

//MAC_2414 replaced by MAC_5827

//MAC_2413 replaced by MAC_5827

//MAC_2412 replaced by MAC_5826

//MAC_2423 replaced by MAC_5827

//MAC_2422 replaced by MAC_5827

//MAC_2421 replaced by MAC_5826

//MAC_2420 replaced by MAC_5827

//MAC_2419 replaced by MAC_5827

//MAC_2418 replaced by MAC_5826

//MAC_2429 replaced by MAC_5827

//MAC_2428 replaced by MAC_5827

//MAC_2427 replaced by MAC_5826

//MAC_2426 replaced by MAC_5827

//MAC_2425 replaced by MAC_5827

//MAC_2424 replaced by MAC_5826

//MAC_2435 replaced by MAC_5827

//MAC_2434 replaced by MAC_5827

//MAC_2433 replaced by MAC_5826

//MAC_2432 replaced by MAC_5827

//MAC_2431 replaced by MAC_5827

//MAC_2430 replaced by MAC_5826

//MAC_2441 replaced by MAC_5827

//MAC_2440 replaced by MAC_5827

//MAC_2439 replaced by MAC_5826

//MAC_2438 replaced by MAC_5827

//MAC_2437 replaced by MAC_5827

//MAC_2436 replaced by MAC_5826

//MAC_2447 replaced by MAC_5827

//MAC_2446 replaced by MAC_5827

//MAC_2445 replaced by MAC_5826

//MAC_2444 replaced by MAC_5827

//MAC_2443 replaced by MAC_5827

//MAC_2442 replaced by MAC_5826

//MAC_2453 replaced by MAC_5827

//MAC_2452 replaced by MAC_5827

//MAC_2451 replaced by MAC_5826

//MAC_2450 replaced by MAC_5827

//MAC_2449 replaced by MAC_5827

//MAC_2448 replaced by MAC_5826

//MAC_2459 replaced by MAC_5827

//MAC_2458 replaced by MAC_5827

//MAC_2457 replaced by MAC_5826

//MAC_2456 replaced by MAC_5827

//MAC_2455 replaced by MAC_5827

//MAC_2454 replaced by MAC_5826

//MAC_2465 replaced by MAC_5827

//MAC_2464 replaced by MAC_5827

//MAC_2463 replaced by MAC_5826

//MAC_2462 replaced by MAC_5827

//MAC_2461 replaced by MAC_5827

//MAC_2460 replaced by MAC_5826

//MAC_2471 replaced by MAC_5827

//MAC_2470 replaced by MAC_5827

//MAC_2469 replaced by MAC_5826

//MAC_2468 replaced by MAC_5827

//MAC_2467 replaced by MAC_5827

//MAC_2466 replaced by MAC_5826

//MAC_2477 replaced by MAC_5827

//MAC_2476 replaced by MAC_5827

//MAC_2475 replaced by MAC_5826

//MAC_2474 replaced by MAC_5827

//MAC_2473 replaced by MAC_5827

//MAC_2472 replaced by MAC_5826

//MAC_2483 replaced by MAC_5827

//MAC_2482 replaced by MAC_5827

//MAC_2481 replaced by MAC_5826

//MAC_2480 replaced by MAC_5827

//MAC_2479 replaced by MAC_5827

//MAC_2478 replaced by MAC_5826

//MAC_2489 replaced by MAC_5827

//MAC_2488 replaced by MAC_5827

//MAC_2487 replaced by MAC_5826

//MAC_2486 replaced by MAC_5827

//MAC_2485 replaced by MAC_5827

//MAC_2484 replaced by MAC_5826

//MAC_2495 replaced by MAC_5827

//MAC_2494 replaced by MAC_5827

//MAC_2493 replaced by MAC_5826

//MAC_2492 replaced by MAC_5827

//MAC_2491 replaced by MAC_5827

//MAC_2490 replaced by MAC_5826

//MAC_2501 replaced by MAC_5827

//MAC_2500 replaced by MAC_5827

//MAC_2499 replaced by MAC_5826

//MAC_2498 replaced by MAC_5827

//MAC_2497 replaced by MAC_5827

//MAC_2496 replaced by MAC_5826

//MAC_2507 replaced by MAC_5827

//MAC_2506 replaced by MAC_5827

//MAC_2505 replaced by MAC_5826

//MAC_2504 replaced by MAC_5827

//MAC_2503 replaced by MAC_5827

//MAC_2502 replaced by MAC_5826

//MAC_2513 replaced by MAC_5827

//MAC_2512 replaced by MAC_5827

//MAC_2511 replaced by MAC_5826

//MAC_2510 replaced by MAC_5827

//MAC_2509 replaced by MAC_5827

//MAC_2508 replaced by MAC_5826

//MAC_2519 replaced by MAC_5827

//MAC_2518 replaced by MAC_5827

//MAC_2517 replaced by MAC_5826

//MAC_2516 replaced by MAC_5827

//MAC_2515 replaced by MAC_5827

//MAC_2514 replaced by MAC_5826

//MAC_2525 replaced by MAC_5827

//MAC_2524 replaced by MAC_5827

//MAC_2523 replaced by MAC_5826

//MAC_2522 replaced by MAC_5827

//MAC_2521 replaced by MAC_5827

//MAC_2520 replaced by MAC_5826

//MAC_2531 replaced by MAC_5827

//MAC_2530 replaced by MAC_5827

//MAC_2529 replaced by MAC_5826

//MAC_2528 replaced by MAC_5827

//MAC_2527 replaced by MAC_5827

//MAC_2526 replaced by MAC_5826

//MAC_2537 replaced by MAC_5827

//MAC_2536 replaced by MAC_5827

//MAC_2535 replaced by MAC_5826

//MAC_2534 replaced by MAC_5827

//MAC_2533 replaced by MAC_5827

//MAC_2532 replaced by MAC_5826

//MAC_2543 replaced by MAC_5827

//MAC_2542 replaced by MAC_5827

//MAC_2541 replaced by MAC_5826

//MAC_2540 replaced by MAC_5827

//MAC_2539 replaced by MAC_5827

//MAC_2538 replaced by MAC_5826

//MAC_2549 replaced by MAC_5827

//MAC_2548 replaced by MAC_5827

//MAC_2547 replaced by MAC_5826

//MAC_2546 replaced by MAC_5827

//MAC_2545 replaced by MAC_5827

//MAC_2544 replaced by MAC_5826

//MAC_2555 replaced by MAC_5827

//MAC_2554 replaced by MAC_5827

//MAC_2553 replaced by MAC_5826

//MAC_2552 replaced by MAC_5827

//MAC_2551 replaced by MAC_5827

//MAC_2550 replaced by MAC_5826

//MAC_2561 replaced by MAC_5827

//MAC_2560 replaced by MAC_5827

//MAC_2559 replaced by MAC_5826

//MAC_2558 replaced by MAC_5827

//MAC_2557 replaced by MAC_5827

//MAC_2556 replaced by MAC_5826

//MAC_2567 replaced by MAC_5827

//MAC_2566 replaced by MAC_5827

//MAC_2565 replaced by MAC_5826

//MAC_2564 replaced by MAC_5827

//MAC_2563 replaced by MAC_5827

//MAC_2562 replaced by MAC_5826

//MAC_2573 replaced by MAC_5827

//MAC_2572 replaced by MAC_5827

//MAC_2571 replaced by MAC_5826

//MAC_2570 replaced by MAC_5827

//MAC_2569 replaced by MAC_5827

//MAC_2568 replaced by MAC_5826

//MAC_2579 replaced by MAC_5827

//MAC_2578 replaced by MAC_5827

//MAC_2577 replaced by MAC_5826

//MAC_2576 replaced by MAC_5827

//MAC_2575 replaced by MAC_5827

//MAC_2574 replaced by MAC_5826

//MAC_2585 replaced by MAC_5827

//MAC_2584 replaced by MAC_5827

//MAC_2583 replaced by MAC_5826

//MAC_2582 replaced by MAC_5827

//MAC_2581 replaced by MAC_5827

//MAC_2580 replaced by MAC_5826

//MAC_2591 replaced by MAC_5827

//MAC_2590 replaced by MAC_5827

//MAC_2589 replaced by MAC_5826

//MAC_2588 replaced by MAC_5827

//MAC_2587 replaced by MAC_5827

//MAC_2586 replaced by MAC_5826

//MAC_2597 replaced by MAC_5827

//MAC_2596 replaced by MAC_5827

//MAC_2595 replaced by MAC_5826

//MAC_2594 replaced by MAC_5827

//MAC_2593 replaced by MAC_5827

//MAC_2592 replaced by MAC_5826

//MAC_2603 replaced by MAC_5827

//MAC_2602 replaced by MAC_5827

//MAC_2601 replaced by MAC_5826

//MAC_2600 replaced by MAC_5827

//MAC_2599 replaced by MAC_5827

//MAC_2598 replaced by MAC_5826

//MAC_2609 replaced by MAC_5827

//MAC_2608 replaced by MAC_5827

//MAC_2607 replaced by MAC_5826

//MAC_2606 replaced by MAC_5827

//MAC_2605 replaced by MAC_5827

//MAC_2604 replaced by MAC_5826

//MAC_2615 replaced by MAC_5827

//MAC_2614 replaced by MAC_5827

//MAC_2613 replaced by MAC_5826

//MAC_2612 replaced by MAC_5827

//MAC_2611 replaced by MAC_5827

//MAC_2610 replaced by MAC_5826

//MAC_2621 replaced by MAC_5827

//MAC_2620 replaced by MAC_5827

//MAC_2619 replaced by MAC_5826

//MAC_2618 replaced by MAC_5827

//MAC_2617 replaced by MAC_5827

//MAC_2616 replaced by MAC_5826

//MAC_2627 replaced by MAC_5827

//MAC_2626 replaced by MAC_5827

//MAC_2625 replaced by MAC_5826

//MAC_2624 replaced by MAC_5827

//MAC_2623 replaced by MAC_5827

//MAC_2622 replaced by MAC_5826

//MAC_2633 replaced by MAC_5827

//MAC_2632 replaced by MAC_5827

//MAC_2631 replaced by MAC_5826

//MAC_2630 replaced by MAC_5827

//MAC_2629 replaced by MAC_5827

//MAC_2628 replaced by MAC_5826

//MAC_2639 replaced by MAC_5827

//MAC_2638 replaced by MAC_5827

//MAC_2637 replaced by MAC_5826

//MAC_2636 replaced by MAC_5827

//MAC_2635 replaced by MAC_5827

//MAC_2634 replaced by MAC_5826

//MAC_2645 replaced by MAC_5827

//MAC_2644 replaced by MAC_5827

//MAC_2643 replaced by MAC_5826

//MAC_2642 replaced by MAC_5827

//MAC_2641 replaced by MAC_5827

//MAC_2640 replaced by MAC_5826

//MAC_2651 replaced by MAC_5827

//MAC_2650 replaced by MAC_5827

//MAC_2649 replaced by MAC_5826

//MAC_2648 replaced by MAC_5827

//MAC_2647 replaced by MAC_5827

//MAC_2646 replaced by MAC_5826

//MAC_2657 replaced by MAC_5827

//MAC_2656 replaced by MAC_5827

//MAC_2655 replaced by MAC_5826

//MAC_2654 replaced by MAC_5827

//MAC_2653 replaced by MAC_5827

//MAC_2652 replaced by MAC_5826

//MAC_2663 replaced by MAC_5827

//MAC_2662 replaced by MAC_5827

//MAC_2661 replaced by MAC_5826

//MAC_2660 replaced by MAC_5827

//MAC_2659 replaced by MAC_5827

//MAC_2658 replaced by MAC_5826

//MAC_2669 replaced by MAC_5827

//MAC_2668 replaced by MAC_5827

//MAC_2667 replaced by MAC_5826

//MAC_2666 replaced by MAC_5827

//MAC_2665 replaced by MAC_5827

//MAC_2664 replaced by MAC_5826

//MAC_2675 replaced by MAC_5827

//MAC_2674 replaced by MAC_5827

//MAC_2673 replaced by MAC_5826

//MAC_2672 replaced by MAC_5827

//MAC_2671 replaced by MAC_5827

//MAC_2670 replaced by MAC_5826

//MAC_2681 replaced by MAC_5827

//MAC_2680 replaced by MAC_5827

//MAC_2679 replaced by MAC_5826

//MAC_2678 replaced by MAC_5827

//MAC_2677 replaced by MAC_5827

//MAC_2676 replaced by MAC_5826

//MAC_2687 replaced by MAC_5827

//MAC_2686 replaced by MAC_5827

//MAC_2685 replaced by MAC_5826

//MAC_2684 replaced by MAC_5827

//MAC_2683 replaced by MAC_5827

//MAC_2682 replaced by MAC_5826

//MAC_2693 replaced by MAC_5827

//MAC_2692 replaced by MAC_5827

//MAC_2691 replaced by MAC_5826

//MAC_2690 replaced by MAC_5827

//MAC_2689 replaced by MAC_5827

//MAC_2688 replaced by MAC_5826

//MAC_2699 replaced by MAC_5827

//MAC_2698 replaced by MAC_5827

//MAC_2697 replaced by MAC_5826

//MAC_2696 replaced by MAC_5827

//MAC_2695 replaced by MAC_5827

//MAC_2694 replaced by MAC_5826

//MAC_2705 replaced by MAC_5827

//MAC_2704 replaced by MAC_5827

//MAC_2703 replaced by MAC_5826

//MAC_2702 replaced by MAC_5827

//MAC_2701 replaced by MAC_5827

//MAC_2700 replaced by MAC_5826

//MAC_2711 replaced by MAC_5827

//MAC_2710 replaced by MAC_5827

//MAC_2709 replaced by MAC_5826

//MAC_2708 replaced by MAC_5827

//MAC_2707 replaced by MAC_5827

//MAC_2706 replaced by MAC_5826

//MAC_2717 replaced by MAC_5827

//MAC_2716 replaced by MAC_5827

//MAC_2715 replaced by MAC_5826

//MAC_2714 replaced by MAC_5827

//MAC_2713 replaced by MAC_5827

//MAC_2712 replaced by MAC_5826

//MAC_2723 replaced by MAC_5827

//MAC_2722 replaced by MAC_5827

//MAC_2721 replaced by MAC_5826

//MAC_2720 replaced by MAC_5827

//MAC_2719 replaced by MAC_5827

//MAC_2718 replaced by MAC_5826

//MAC_2729 replaced by MAC_5827

//MAC_2728 replaced by MAC_5827

//MAC_2727 replaced by MAC_5826

//MAC_2726 replaced by MAC_5827

//MAC_2725 replaced by MAC_5827

//MAC_2724 replaced by MAC_5826

//MAC_2735 replaced by MAC_5827

//MAC_2734 replaced by MAC_5827

//MAC_2733 replaced by MAC_5826

//MAC_2732 replaced by MAC_5827

//MAC_2731 replaced by MAC_5827

//MAC_2730 replaced by MAC_5826

//MAC_2741 replaced by MAC_5827

//MAC_2740 replaced by MAC_5827

//MAC_2739 replaced by MAC_5826

//MAC_2738 replaced by MAC_5827

//MAC_2737 replaced by MAC_5827

//MAC_2736 replaced by MAC_5826

//MAC_2747 replaced by MAC_5827

//MAC_2746 replaced by MAC_5827

//MAC_2745 replaced by MAC_5826

//MAC_2744 replaced by MAC_5827

//MAC_2743 replaced by MAC_5827

//MAC_2742 replaced by MAC_5826

//MAC_2753 replaced by MAC_5827

//MAC_2752 replaced by MAC_5827

//MAC_2751 replaced by MAC_5826

//MAC_2750 replaced by MAC_5827

//MAC_2749 replaced by MAC_5827

//MAC_2748 replaced by MAC_5826

//MAC_2759 replaced by MAC_5827

//MAC_2758 replaced by MAC_5827

//MAC_2757 replaced by MAC_5826

//MAC_2756 replaced by MAC_5827

//MAC_2755 replaced by MAC_5827

//MAC_2754 replaced by MAC_5826

//MAC_2765 replaced by MAC_5827

//MAC_2764 replaced by MAC_5827

//MAC_2763 replaced by MAC_5826

//MAC_2762 replaced by MAC_5827

//MAC_2761 replaced by MAC_5827

//MAC_2760 replaced by MAC_5826

//MAC_2771 replaced by MAC_5827

//MAC_2770 replaced by MAC_5827

//MAC_2769 replaced by MAC_5826

//MAC_2768 replaced by MAC_5827

//MAC_2767 replaced by MAC_5827

//MAC_2766 replaced by MAC_5826

//MAC_2777 replaced by MAC_5827

//MAC_2776 replaced by MAC_5827

//MAC_2775 replaced by MAC_5826

//MAC_2774 replaced by MAC_5827

//MAC_2773 replaced by MAC_5827

//MAC_2772 replaced by MAC_5826

//MAC_2783 replaced by MAC_5827

//MAC_2782 replaced by MAC_5827

//MAC_2781 replaced by MAC_5826

//MAC_2780 replaced by MAC_5827

//MAC_2779 replaced by MAC_5827

//MAC_2778 replaced by MAC_5826

//MAC_2789 replaced by MAC_5827

//MAC_2788 replaced by MAC_5827

//MAC_2787 replaced by MAC_5826

//MAC_2786 replaced by MAC_5827

//MAC_2785 replaced by MAC_5827

//MAC_2784 replaced by MAC_5826

//MAC_2795 replaced by MAC_5827

//MAC_2794 replaced by MAC_5827

//MAC_2793 replaced by MAC_5826

//MAC_2792 replaced by MAC_5827

//MAC_2791 replaced by MAC_5827

//MAC_2790 replaced by MAC_5826

//MAC_2801 replaced by MAC_5827

//MAC_2800 replaced by MAC_5827

//MAC_2799 replaced by MAC_5826

//MAC_2798 replaced by MAC_5827

//MAC_2797 replaced by MAC_5827

//MAC_2796 replaced by MAC_5826

//MAC_2807 replaced by MAC_5827

//MAC_2806 replaced by MAC_5827

//MAC_2805 replaced by MAC_5826

//MAC_2804 replaced by MAC_5827

//MAC_2803 replaced by MAC_5827

//MAC_2802 replaced by MAC_5826

//MAC_2813 replaced by MAC_5827

//MAC_2812 replaced by MAC_5827

//MAC_2811 replaced by MAC_5826

//MAC_2810 replaced by MAC_5827

//MAC_2809 replaced by MAC_5827

//MAC_2808 replaced by MAC_5826

//MAC_2819 replaced by MAC_5827

//MAC_2818 replaced by MAC_5827

//MAC_2817 replaced by MAC_5826

//MAC_2816 replaced by MAC_5827

//MAC_2815 replaced by MAC_5827

//MAC_2814 replaced by MAC_5826

//MAC_2825 replaced by MAC_5827

//MAC_2824 replaced by MAC_5827

//MAC_2823 replaced by MAC_5826

//MAC_2822 replaced by MAC_5827

//MAC_2821 replaced by MAC_5827

//MAC_2820 replaced by MAC_5826

//MAC_2831 replaced by MAC_5827

//MAC_2830 replaced by MAC_5827

//MAC_2829 replaced by MAC_5826

//MAC_2828 replaced by MAC_5827

//MAC_2827 replaced by MAC_5827

//MAC_2826 replaced by MAC_5826

//MAC_2837 replaced by MAC_5827

//MAC_2836 replaced by MAC_5827

//MAC_2835 replaced by MAC_5826

//MAC_2834 replaced by MAC_5827

//MAC_2833 replaced by MAC_5827

//MAC_2832 replaced by MAC_5826

//MAC_2843 replaced by MAC_5827

//MAC_2842 replaced by MAC_5827

//MAC_2841 replaced by MAC_5826

//MAC_2840 replaced by MAC_5827

//MAC_2839 replaced by MAC_5827

//MAC_2838 replaced by MAC_5826

//MAC_2849 replaced by MAC_5827

//MAC_2848 replaced by MAC_5827

//MAC_2847 replaced by MAC_5826

//MAC_2846 replaced by MAC_5827

//MAC_2845 replaced by MAC_5827

//MAC_2844 replaced by MAC_5826

//MAC_2855 replaced by MAC_5827

//MAC_2854 replaced by MAC_5827

//MAC_2853 replaced by MAC_5826

//MAC_2852 replaced by MAC_5827

//MAC_2851 replaced by MAC_5827

//MAC_2850 replaced by MAC_5826

//MAC_2861 replaced by MAC_5827

//MAC_2860 replaced by MAC_5827

//MAC_2859 replaced by MAC_5826

//MAC_2858 replaced by MAC_5827

//MAC_2857 replaced by MAC_5827

//MAC_2856 replaced by MAC_5826

//MAC_2867 replaced by MAC_5827

//MAC_2866 replaced by MAC_5827

//MAC_2865 replaced by MAC_5826

//MAC_2864 replaced by MAC_5827

//MAC_2863 replaced by MAC_5827

//MAC_2862 replaced by MAC_5826

//MAC_2873 replaced by MAC_5827

//MAC_2872 replaced by MAC_5827

//MAC_2871 replaced by MAC_5826

//MAC_2870 replaced by MAC_5827

//MAC_2869 replaced by MAC_5827

//MAC_2868 replaced by MAC_5826

//MAC_2879 replaced by MAC_5827

//MAC_2878 replaced by MAC_5827

//MAC_2877 replaced by MAC_5826

//MAC_2876 replaced by MAC_5827

//MAC_2875 replaced by MAC_5827

//MAC_2874 replaced by MAC_5826

//MAC_2885 replaced by MAC_5827

//MAC_2884 replaced by MAC_5827

//MAC_2883 replaced by MAC_5826

//MAC_2882 replaced by MAC_5827

//MAC_2881 replaced by MAC_5827

//MAC_2880 replaced by MAC_5826

//MAC_2891 replaced by MAC_5827

//MAC_2890 replaced by MAC_5827

//MAC_2889 replaced by MAC_5826

//MAC_2888 replaced by MAC_5827

//MAC_2887 replaced by MAC_5827

//MAC_2886 replaced by MAC_5826

//MAC_2897 replaced by MAC_5827

//MAC_2896 replaced by MAC_5827

//MAC_2895 replaced by MAC_5826

//MAC_2894 replaced by MAC_5827

//MAC_2893 replaced by MAC_5827

//MAC_2892 replaced by MAC_5826

//MAC_2903 replaced by MAC_5827

//MAC_2902 replaced by MAC_5827

//MAC_2901 replaced by MAC_5826

//MAC_2900 replaced by MAC_5827

//MAC_2899 replaced by MAC_5827

//MAC_2898 replaced by MAC_5826

//MAC_2909 replaced by MAC_5827

//MAC_2908 replaced by MAC_5827

//MAC_2907 replaced by MAC_5826

//MAC_2906 replaced by MAC_5827

//MAC_2905 replaced by MAC_5827

//MAC_2904 replaced by MAC_5826

//MAC_2915 replaced by MAC_5827

//MAC_2914 replaced by MAC_5827

//MAC_2913 replaced by MAC_5826

//MAC_2912 replaced by MAC_5827

//MAC_2911 replaced by MAC_5827

//MAC_2910 replaced by MAC_5826

//MAC_2921 replaced by MAC_5827

//MAC_2920 replaced by MAC_5827

//MAC_2919 replaced by MAC_5826

//MAC_2918 replaced by MAC_5827

//MAC_2917 replaced by MAC_5827

//MAC_2916 replaced by MAC_5826

//MAC_2927 replaced by MAC_5827

//MAC_2926 replaced by MAC_5827

//MAC_2925 replaced by MAC_5826

//MAC_2924 replaced by MAC_5827

//MAC_2923 replaced by MAC_5827

//MAC_2922 replaced by MAC_5826

//MAC_2933 replaced by MAC_5827

//MAC_2932 replaced by MAC_5827

//MAC_2931 replaced by MAC_5826

//MAC_2930 replaced by MAC_5827

//MAC_2929 replaced by MAC_5827

//MAC_2928 replaced by MAC_5826

//MAC_2939 replaced by MAC_5827

//MAC_2938 replaced by MAC_5827

//MAC_2937 replaced by MAC_5826

//MAC_2936 replaced by MAC_5827

//MAC_2935 replaced by MAC_5827

//MAC_2934 replaced by MAC_5826

//MAC_2945 replaced by MAC_5827

//MAC_2944 replaced by MAC_5827

//MAC_2943 replaced by MAC_5826

//MAC_2942 replaced by MAC_5827

//MAC_2941 replaced by MAC_5827

//MAC_2940 replaced by MAC_5826

//MAC_2951 replaced by MAC_5827

//MAC_2950 replaced by MAC_5827

//MAC_2949 replaced by MAC_5826

//MAC_2948 replaced by MAC_5827

//MAC_2947 replaced by MAC_5827

//MAC_2946 replaced by MAC_5826

//MAC_2957 replaced by MAC_5827

//MAC_2956 replaced by MAC_5827

//MAC_2955 replaced by MAC_5826

//MAC_2954 replaced by MAC_5827

//MAC_2953 replaced by MAC_5827

//MAC_2952 replaced by MAC_5826

//MAC_2963 replaced by MAC_5827

//MAC_2962 replaced by MAC_5827

//MAC_2961 replaced by MAC_5826

//MAC_2960 replaced by MAC_5827

//MAC_2959 replaced by MAC_5827

//MAC_2958 replaced by MAC_5826

//MAC_2969 replaced by MAC_5827

//MAC_2968 replaced by MAC_5827

//MAC_2967 replaced by MAC_5826

//MAC_2966 replaced by MAC_5827

//MAC_2965 replaced by MAC_5827

//MAC_2964 replaced by MAC_5826

//MAC_2975 replaced by MAC_5827

//MAC_2974 replaced by MAC_5827

//MAC_2973 replaced by MAC_5826

//MAC_2972 replaced by MAC_5827

//MAC_2971 replaced by MAC_5827

//MAC_2970 replaced by MAC_5826

//MAC_2981 replaced by MAC_5827

//MAC_2980 replaced by MAC_5827

//MAC_2979 replaced by MAC_5826

//MAC_2978 replaced by MAC_5827

//MAC_2977 replaced by MAC_5827

//MAC_2976 replaced by MAC_5826

//MAC_2987 replaced by MAC_5827

//MAC_2986 replaced by MAC_5827

//MAC_2985 replaced by MAC_5826

//MAC_2984 replaced by MAC_5827

//MAC_2983 replaced by MAC_5827

//MAC_2982 replaced by MAC_5826

//MAC_2993 replaced by MAC_5827

//MAC_2992 replaced by MAC_5827

//MAC_2991 replaced by MAC_5826

//MAC_2990 replaced by MAC_5827

//MAC_2989 replaced by MAC_5827

//MAC_2988 replaced by MAC_5826

//MAC_2999 replaced by MAC_5827

//MAC_2998 replaced by MAC_5827

//MAC_2997 replaced by MAC_5826

//MAC_2996 replaced by MAC_5827

//MAC_2995 replaced by MAC_5827

//MAC_2994 replaced by MAC_5826

//MAC_3005 replaced by MAC_5827

//MAC_3004 replaced by MAC_5827

//MAC_3003 replaced by MAC_5826

//MAC_3002 replaced by MAC_5827

//MAC_3001 replaced by MAC_5827

//MAC_3000 replaced by MAC_5826

//MAC_3011 replaced by MAC_5827

//MAC_3010 replaced by MAC_5827

//MAC_3009 replaced by MAC_5826

//MAC_3008 replaced by MAC_5827

//MAC_3007 replaced by MAC_5827

//MAC_3006 replaced by MAC_5826

//MAC_3017 replaced by MAC_5827

//MAC_3016 replaced by MAC_5827

//MAC_3015 replaced by MAC_5826

//MAC_3014 replaced by MAC_5827

//MAC_3013 replaced by MAC_5827

//MAC_3012 replaced by MAC_5826

//MAC_3023 replaced by MAC_5827

//MAC_3022 replaced by MAC_5827

//MAC_3021 replaced by MAC_5826

//MAC_3020 replaced by MAC_5827

//MAC_3019 replaced by MAC_5827

//MAC_3018 replaced by MAC_5826

//MAC_3029 replaced by MAC_5827

//MAC_3028 replaced by MAC_5827

//MAC_3027 replaced by MAC_5826

//MAC_3026 replaced by MAC_5827

//MAC_3025 replaced by MAC_5827

//MAC_3024 replaced by MAC_5826

//MAC_3035 replaced by MAC_5827

//MAC_3034 replaced by MAC_5827

//MAC_3033 replaced by MAC_5826

//MAC_3032 replaced by MAC_5827

//MAC_3031 replaced by MAC_5827

//MAC_3030 replaced by MAC_5826

//MAC_3041 replaced by MAC_5827

//MAC_3040 replaced by MAC_5827

//MAC_3039 replaced by MAC_5826

//MAC_3038 replaced by MAC_5827

//MAC_3037 replaced by MAC_5827

//MAC_3036 replaced by MAC_5826

//MAC_3047 replaced by MAC_5827

//MAC_3046 replaced by MAC_5827

//MAC_3045 replaced by MAC_5826

//MAC_3044 replaced by MAC_5827

//MAC_3043 replaced by MAC_5827

//MAC_3042 replaced by MAC_5826

//MAC_3053 replaced by MAC_5827

//MAC_3052 replaced by MAC_5827

//MAC_3051 replaced by MAC_5826

//MAC_3050 replaced by MAC_5827

//MAC_3049 replaced by MAC_5827

//MAC_3048 replaced by MAC_5826

//MAC_3059 replaced by MAC_5827

//MAC_3058 replaced by MAC_5827

//MAC_3057 replaced by MAC_5826

//MAC_3056 replaced by MAC_5827

//MAC_3055 replaced by MAC_5827

//MAC_3054 replaced by MAC_5826

//MAC_3065 replaced by MAC_5827

//MAC_3064 replaced by MAC_5827

//MAC_3063 replaced by MAC_5826

//MAC_3062 replaced by MAC_5827

//MAC_3061 replaced by MAC_5827

//MAC_3060 replaced by MAC_5826

//MAC_3071 replaced by MAC_5827

//MAC_3070 replaced by MAC_5827

//MAC_3069 replaced by MAC_5826

//MAC_3068 replaced by MAC_5827

//MAC_3067 replaced by MAC_5827

//MAC_3066 replaced by MAC_5826

//MAC_3077 replaced by MAC_5827

//MAC_3076 replaced by MAC_5827

//MAC_3075 replaced by MAC_5826

//MAC_3074 replaced by MAC_5827

//MAC_3073 replaced by MAC_5827

//MAC_3072 replaced by MAC_5826

//MAC_3083 replaced by MAC_5827

//MAC_3082 replaced by MAC_5827

//MAC_3081 replaced by MAC_5826

//MAC_3080 replaced by MAC_5827

//MAC_3079 replaced by MAC_5827

//MAC_3078 replaced by MAC_5826

//MAC_3089 replaced by MAC_5827

//MAC_3088 replaced by MAC_5827

//MAC_3087 replaced by MAC_5826

//MAC_3086 replaced by MAC_5827

//MAC_3085 replaced by MAC_5827

//MAC_3084 replaced by MAC_5826

//MAC_3095 replaced by MAC_5827

//MAC_3094 replaced by MAC_5827

//MAC_3093 replaced by MAC_5826

//MAC_3092 replaced by MAC_5827

//MAC_3091 replaced by MAC_5827

//MAC_3090 replaced by MAC_5826

//MAC_3101 replaced by MAC_5827

//MAC_3100 replaced by MAC_5827

//MAC_3099 replaced by MAC_5826

//MAC_3098 replaced by MAC_5827

//MAC_3097 replaced by MAC_5827

//MAC_3096 replaced by MAC_5826

//MAC_3107 replaced by MAC_5827

//MAC_3106 replaced by MAC_5827

//MAC_3105 replaced by MAC_5826

//MAC_3104 replaced by MAC_5827

//MAC_3103 replaced by MAC_5827

//MAC_3102 replaced by MAC_5826

//MAC_3113 replaced by MAC_5827

//MAC_3112 replaced by MAC_5827

//MAC_3111 replaced by MAC_5826

//MAC_3110 replaced by MAC_5827

//MAC_3109 replaced by MAC_5827

//MAC_3108 replaced by MAC_5826

//MAC_3119 replaced by MAC_5827

//MAC_3118 replaced by MAC_5827

//MAC_3117 replaced by MAC_5826

//MAC_3116 replaced by MAC_5827

//MAC_3115 replaced by MAC_5827

//MAC_3114 replaced by MAC_5826

//MAC_3125 replaced by MAC_5827

//MAC_3124 replaced by MAC_5827

//MAC_3123 replaced by MAC_5826

//MAC_3122 replaced by MAC_5827

//MAC_3121 replaced by MAC_5827

//MAC_3120 replaced by MAC_5826

//MAC_3131 replaced by MAC_5827

//MAC_3130 replaced by MAC_5827

//MAC_3129 replaced by MAC_5826

//MAC_3128 replaced by MAC_5827

//MAC_3127 replaced by MAC_5827

//MAC_3126 replaced by MAC_5826

//MAC_3137 replaced by MAC_5827

//MAC_3136 replaced by MAC_5827

//MAC_3135 replaced by MAC_5826

//MAC_3134 replaced by MAC_5827

//MAC_3133 replaced by MAC_5827

//MAC_3132 replaced by MAC_5826

//MAC_3143 replaced by MAC_5827

//MAC_3142 replaced by MAC_5827

//MAC_3141 replaced by MAC_5826

//MAC_3140 replaced by MAC_5827

//MAC_3139 replaced by MAC_5827

//MAC_3138 replaced by MAC_5826

//MAC_3149 replaced by MAC_5827

//MAC_3148 replaced by MAC_5827

//MAC_3147 replaced by MAC_5826

//MAC_3146 replaced by MAC_5827

//MAC_3145 replaced by MAC_5827

//MAC_3144 replaced by MAC_5826

//MAC_3155 replaced by MAC_5827

//MAC_3154 replaced by MAC_5827

//MAC_3153 replaced by MAC_5826

//MAC_3152 replaced by MAC_5827

//MAC_3151 replaced by MAC_5827

//MAC_3150 replaced by MAC_5826

//MAC_3161 replaced by MAC_5827

//MAC_3160 replaced by MAC_5827

//MAC_3159 replaced by MAC_5826

//MAC_3158 replaced by MAC_5827

//MAC_3157 replaced by MAC_5827

//MAC_3156 replaced by MAC_5826

//MAC_3167 replaced by MAC_5827

//MAC_3166 replaced by MAC_5827

//MAC_3165 replaced by MAC_5826

//MAC_3164 replaced by MAC_5827

//MAC_3163 replaced by MAC_5827

//MAC_3162 replaced by MAC_5826

//MAC_3173 replaced by MAC_5827

//MAC_3172 replaced by MAC_5827

//MAC_3171 replaced by MAC_5826

//MAC_3170 replaced by MAC_5827

//MAC_3169 replaced by MAC_5827

//MAC_3168 replaced by MAC_5826

//MAC_3179 replaced by MAC_5827

//MAC_3178 replaced by MAC_5827

//MAC_3177 replaced by MAC_5826

//MAC_3176 replaced by MAC_5827

//MAC_3175 replaced by MAC_5827

//MAC_3174 replaced by MAC_5826

//MAC_3185 replaced by MAC_5827

//MAC_3184 replaced by MAC_5827

//MAC_3183 replaced by MAC_5826

//MAC_3182 replaced by MAC_5827

//MAC_3181 replaced by MAC_5827

//MAC_3180 replaced by MAC_5826

//MAC_3191 replaced by MAC_5827

//MAC_3190 replaced by MAC_5827

//MAC_3189 replaced by MAC_5826

//MAC_3188 replaced by MAC_5827

//MAC_3187 replaced by MAC_5827

//MAC_3186 replaced by MAC_5826

//MAC_3197 replaced by MAC_5827

//MAC_3196 replaced by MAC_5827

//MAC_3195 replaced by MAC_5826

//MAC_3194 replaced by MAC_5827

//MAC_3193 replaced by MAC_5827

//MAC_3192 replaced by MAC_5826

//MAC_3203 replaced by MAC_5827

//MAC_3202 replaced by MAC_5827

//MAC_3201 replaced by MAC_5826

//MAC_3200 replaced by MAC_5827

//MAC_3199 replaced by MAC_5827

//MAC_3198 replaced by MAC_5826

//MAC_3209 replaced by MAC_5827

//MAC_3208 replaced by MAC_5827

//MAC_3207 replaced by MAC_5826

//MAC_3206 replaced by MAC_5827

//MAC_3205 replaced by MAC_5827

//MAC_3204 replaced by MAC_5826

//MAC_3215 replaced by MAC_5827

//MAC_3214 replaced by MAC_5827

//MAC_3213 replaced by MAC_5826

//MAC_3212 replaced by MAC_5827

//MAC_3211 replaced by MAC_5827

//MAC_3210 replaced by MAC_5826

//MAC_3221 replaced by MAC_5827

//MAC_3220 replaced by MAC_5827

//MAC_3219 replaced by MAC_5826

//MAC_3218 replaced by MAC_5827

//MAC_3217 replaced by MAC_5827

//MAC_3216 replaced by MAC_5826

//MAC_3227 replaced by MAC_5827

//MAC_3226 replaced by MAC_5827

//MAC_3225 replaced by MAC_5826

//MAC_3224 replaced by MAC_5827

//MAC_3223 replaced by MAC_5827

//MAC_3222 replaced by MAC_5826

//MAC_3233 replaced by MAC_5827

//MAC_3232 replaced by MAC_5827

//MAC_3231 replaced by MAC_5826

//MAC_3230 replaced by MAC_5827

//MAC_3229 replaced by MAC_5827

//MAC_3228 replaced by MAC_5826

//MAC_3239 replaced by MAC_5827

//MAC_3238 replaced by MAC_5827

//MAC_3237 replaced by MAC_5826

//MAC_3236 replaced by MAC_5827

//MAC_3235 replaced by MAC_5827

//MAC_3234 replaced by MAC_5826

//MAC_3245 replaced by MAC_5827

//MAC_3244 replaced by MAC_5827

//MAC_3243 replaced by MAC_5826

//MAC_3242 replaced by MAC_5827

//MAC_3241 replaced by MAC_5827

//MAC_3240 replaced by MAC_5826

//MAC_3251 replaced by MAC_5827

//MAC_3250 replaced by MAC_5827

//MAC_3249 replaced by MAC_5826

//MAC_3248 replaced by MAC_5827

//MAC_3247 replaced by MAC_5827

//MAC_3246 replaced by MAC_5826

//MAC_3257 replaced by MAC_5827

//MAC_3256 replaced by MAC_5827

//MAC_3255 replaced by MAC_5826

//MAC_3254 replaced by MAC_5827

//MAC_3253 replaced by MAC_5827

//MAC_3252 replaced by MAC_5826

//MAC_3263 replaced by MAC_5827

//MAC_3262 replaced by MAC_5827

//MAC_3261 replaced by MAC_5826

//MAC_3260 replaced by MAC_5827

//MAC_3259 replaced by MAC_5827

//MAC_3258 replaced by MAC_5826

//MAC_3269 replaced by MAC_5827

//MAC_3268 replaced by MAC_5827

//MAC_3267 replaced by MAC_5826

//MAC_3266 replaced by MAC_5827

//MAC_3265 replaced by MAC_5827

//MAC_3264 replaced by MAC_5826

//MAC_3275 replaced by MAC_5827

//MAC_3274 replaced by MAC_5827

//MAC_3273 replaced by MAC_5826

//MAC_3272 replaced by MAC_5827

//MAC_3271 replaced by MAC_5827

//MAC_3270 replaced by MAC_5826

//MAC_3281 replaced by MAC_5827

//MAC_3280 replaced by MAC_5827

//MAC_3279 replaced by MAC_5826

//MAC_3278 replaced by MAC_5827

//MAC_3277 replaced by MAC_5827

//MAC_3276 replaced by MAC_5826

//MAC_3287 replaced by MAC_5827

//MAC_3286 replaced by MAC_5827

//MAC_3285 replaced by MAC_5826

//MAC_3284 replaced by MAC_5827

//MAC_3283 replaced by MAC_5827

//MAC_3282 replaced by MAC_5826

//MAC_3293 replaced by MAC_5827

//MAC_3292 replaced by MAC_5827

//MAC_3291 replaced by MAC_5826

//MAC_3290 replaced by MAC_5827

//MAC_3289 replaced by MAC_5827

//MAC_3288 replaced by MAC_5826

//MAC_3299 replaced by MAC_5827

//MAC_3298 replaced by MAC_5827

//MAC_3297 replaced by MAC_5826

//MAC_3296 replaced by MAC_5827

//MAC_3295 replaced by MAC_5827

//MAC_3294 replaced by MAC_5826

//MAC_3305 replaced by MAC_5827

//MAC_3304 replaced by MAC_5827

//MAC_3303 replaced by MAC_5826

//MAC_3302 replaced by MAC_5827

//MAC_3301 replaced by MAC_5827

//MAC_3300 replaced by MAC_5826

//MAC_3311 replaced by MAC_5827

//MAC_3310 replaced by MAC_5827

//MAC_3309 replaced by MAC_5826

//MAC_3308 replaced by MAC_5827

//MAC_3307 replaced by MAC_5827

//MAC_3306 replaced by MAC_5826

//MAC_3317 replaced by MAC_5827

//MAC_3316 replaced by MAC_5827

//MAC_3315 replaced by MAC_5826

//MAC_3314 replaced by MAC_5827

//MAC_3313 replaced by MAC_5827

//MAC_3312 replaced by MAC_5826

//MAC_3323 replaced by MAC_5827

//MAC_3322 replaced by MAC_5827

//MAC_3321 replaced by MAC_5826

//MAC_3320 replaced by MAC_5827

//MAC_3319 replaced by MAC_5827

//MAC_3318 replaced by MAC_5826

//MAC_3329 replaced by MAC_5827

//MAC_3328 replaced by MAC_5827

//MAC_3327 replaced by MAC_5826

//MAC_3326 replaced by MAC_5827

//MAC_3325 replaced by MAC_5827

//MAC_3324 replaced by MAC_5826

//MAC_3335 replaced by MAC_5827

//MAC_3334 replaced by MAC_5827

//MAC_3333 replaced by MAC_5826

//MAC_3332 replaced by MAC_5827

//MAC_3331 replaced by MAC_5827

//MAC_3330 replaced by MAC_5826

//MAC_3341 replaced by MAC_5827

//MAC_3340 replaced by MAC_5827

//MAC_3339 replaced by MAC_5826

//MAC_3338 replaced by MAC_5827

//MAC_3337 replaced by MAC_5827

//MAC_3336 replaced by MAC_5826

//MAC_3347 replaced by MAC_5827

//MAC_3346 replaced by MAC_5827

//MAC_3345 replaced by MAC_5826

//MAC_3344 replaced by MAC_5827

//MAC_3343 replaced by MAC_5827

//MAC_3342 replaced by MAC_5826

//MAC_3353 replaced by MAC_5827

//MAC_3352 replaced by MAC_5827

//MAC_3351 replaced by MAC_5826

//MAC_3350 replaced by MAC_5827

//MAC_3349 replaced by MAC_5827

//MAC_3348 replaced by MAC_5826

//MAC_3359 replaced by MAC_5827

//MAC_3358 replaced by MAC_5827

//MAC_3357 replaced by MAC_5826

//MAC_3356 replaced by MAC_5827

//MAC_3355 replaced by MAC_5827

//MAC_3354 replaced by MAC_5826

//MAC_3365 replaced by MAC_5827

//MAC_3364 replaced by MAC_5827

//MAC_3363 replaced by MAC_5826

//MAC_3362 replaced by MAC_5827

//MAC_3361 replaced by MAC_5827

//MAC_3360 replaced by MAC_5826

//MAC_3371 replaced by MAC_5827

//MAC_3370 replaced by MAC_5827

//MAC_3369 replaced by MAC_5826

//MAC_3368 replaced by MAC_5827

//MAC_3367 replaced by MAC_5827

//MAC_3366 replaced by MAC_5826

//MAC_3377 replaced by MAC_5827

//MAC_3376 replaced by MAC_5827

//MAC_3375 replaced by MAC_5826

//MAC_3374 replaced by MAC_5827

//MAC_3373 replaced by MAC_5827

//MAC_3372 replaced by MAC_5826

//MAC_3383 replaced by MAC_5827

//MAC_3382 replaced by MAC_5827

//MAC_3381 replaced by MAC_5826

//MAC_3380 replaced by MAC_5827

//MAC_3379 replaced by MAC_5827

//MAC_3378 replaced by MAC_5826

//MAC_3389 replaced by MAC_5827

//MAC_3388 replaced by MAC_5827

//MAC_3387 replaced by MAC_5826

//MAC_3386 replaced by MAC_5827

//MAC_3385 replaced by MAC_5827

//MAC_3384 replaced by MAC_5826

//MAC_3395 replaced by MAC_5827

//MAC_3394 replaced by MAC_5827

//MAC_3393 replaced by MAC_5826

//MAC_3392 replaced by MAC_5827

//MAC_3391 replaced by MAC_5827

//MAC_3390 replaced by MAC_5826

//MAC_3401 replaced by MAC_5827

//MAC_3400 replaced by MAC_5827

//MAC_3399 replaced by MAC_5826

//MAC_3398 replaced by MAC_5827

//MAC_3397 replaced by MAC_5827

//MAC_3396 replaced by MAC_5826

//MAC_3407 replaced by MAC_5827

//MAC_3406 replaced by MAC_5827

//MAC_3405 replaced by MAC_5826

//MAC_3404 replaced by MAC_5827

//MAC_3403 replaced by MAC_5827

//MAC_3402 replaced by MAC_5826

//MAC_3413 replaced by MAC_5827

//MAC_3412 replaced by MAC_5827

//MAC_3411 replaced by MAC_5826

//MAC_3410 replaced by MAC_5827

//MAC_3409 replaced by MAC_5827

//MAC_3408 replaced by MAC_5826

//MAC_3419 replaced by MAC_5827

//MAC_3418 replaced by MAC_5827

//MAC_3417 replaced by MAC_5826

//MAC_3416 replaced by MAC_5827

//MAC_3415 replaced by MAC_5827

//MAC_3414 replaced by MAC_5826

//MAC_3425 replaced by MAC_5827

//MAC_3424 replaced by MAC_5827

//MAC_3423 replaced by MAC_5826

//MAC_3422 replaced by MAC_5827

//MAC_3421 replaced by MAC_5827

//MAC_3420 replaced by MAC_5826

//MAC_3431 replaced by MAC_5827

//MAC_3430 replaced by MAC_5827

//MAC_3429 replaced by MAC_5826

//MAC_3428 replaced by MAC_5827

//MAC_3427 replaced by MAC_5827

//MAC_3426 replaced by MAC_5826

//MAC_3437 replaced by MAC_5827

//MAC_3436 replaced by MAC_5827

//MAC_3435 replaced by MAC_5826

//MAC_3434 replaced by MAC_5827

//MAC_3433 replaced by MAC_5827

//MAC_3432 replaced by MAC_5826

//MAC_3443 replaced by MAC_5827

//MAC_3442 replaced by MAC_5827

//MAC_3441 replaced by MAC_5826

//MAC_3440 replaced by MAC_5827

//MAC_3439 replaced by MAC_5827

//MAC_3438 replaced by MAC_5826

//MAC_3449 replaced by MAC_5827

//MAC_3448 replaced by MAC_5827

//MAC_3447 replaced by MAC_5826

//MAC_3446 replaced by MAC_5827

//MAC_3445 replaced by MAC_5827

//MAC_3444 replaced by MAC_5826

//MAC_3455 replaced by MAC_5827

//MAC_3454 replaced by MAC_5827

//MAC_3453 replaced by MAC_5826

//MAC_3452 replaced by MAC_5827

//MAC_3451 replaced by MAC_5827

//MAC_3450 replaced by MAC_5826

//MAC_3461 replaced by MAC_5827

//MAC_3460 replaced by MAC_5827

//MAC_3459 replaced by MAC_5826

//MAC_3458 replaced by MAC_5827

//MAC_3457 replaced by MAC_5827

//MAC_3456 replaced by MAC_5826

//MAC_3467 replaced by MAC_5827

//MAC_3466 replaced by MAC_5827

//MAC_3465 replaced by MAC_5826

//MAC_3464 replaced by MAC_5827

//MAC_3463 replaced by MAC_5827

//MAC_3462 replaced by MAC_5826

//MAC_3473 replaced by MAC_5827

//MAC_3472 replaced by MAC_5827

//MAC_3471 replaced by MAC_5826

//MAC_3470 replaced by MAC_5827

//MAC_3469 replaced by MAC_5827

//MAC_3468 replaced by MAC_5826

//MAC_3479 replaced by MAC_5827

//MAC_3478 replaced by MAC_5827

//MAC_3477 replaced by MAC_5826

//MAC_3476 replaced by MAC_5827

//MAC_3475 replaced by MAC_5827

//MAC_3474 replaced by MAC_5826

//MAC_3485 replaced by MAC_5827

//MAC_3484 replaced by MAC_5827

//MAC_3483 replaced by MAC_5826

//MAC_3482 replaced by MAC_5827

//MAC_3481 replaced by MAC_5827

//MAC_3480 replaced by MAC_5826

//MAC_3491 replaced by MAC_5827

//MAC_3490 replaced by MAC_5827

//MAC_3489 replaced by MAC_5826

//MAC_3488 replaced by MAC_5827

//MAC_3487 replaced by MAC_5827

//MAC_3486 replaced by MAC_5826

//MAC_3497 replaced by MAC_5827

//MAC_3496 replaced by MAC_5827

//MAC_3495 replaced by MAC_5826

//MAC_3494 replaced by MAC_5827

//MAC_3493 replaced by MAC_5827

//MAC_3492 replaced by MAC_5826

//MAC_3503 replaced by MAC_5827

//MAC_3502 replaced by MAC_5827

//MAC_3501 replaced by MAC_5826

//MAC_3500 replaced by MAC_5827

//MAC_3499 replaced by MAC_5827

//MAC_3498 replaced by MAC_5826

//MAC_3509 replaced by MAC_5827

//MAC_3508 replaced by MAC_5827

//MAC_3507 replaced by MAC_5826

//MAC_3506 replaced by MAC_5827

//MAC_3505 replaced by MAC_5827

//MAC_3504 replaced by MAC_5826

//MAC_3515 replaced by MAC_5827

//MAC_3514 replaced by MAC_5827

//MAC_3513 replaced by MAC_5826

//MAC_3512 replaced by MAC_5827

//MAC_3511 replaced by MAC_5827

//MAC_3510 replaced by MAC_5826

//MAC_3521 replaced by MAC_5827

//MAC_3520 replaced by MAC_5827

//MAC_3519 replaced by MAC_5826

//MAC_3518 replaced by MAC_5827

//MAC_3517 replaced by MAC_5827

//MAC_3516 replaced by MAC_5826

//MAC_3527 replaced by MAC_5827

//MAC_3526 replaced by MAC_5827

//MAC_3525 replaced by MAC_5826

//MAC_3524 replaced by MAC_5827

//MAC_3523 replaced by MAC_5827

//MAC_3522 replaced by MAC_5826

//MAC_3533 replaced by MAC_5827

//MAC_3532 replaced by MAC_5827

//MAC_3531 replaced by MAC_5826

//MAC_3530 replaced by MAC_5827

//MAC_3529 replaced by MAC_5827

//MAC_3528 replaced by MAC_5826

//MAC_3539 replaced by MAC_5827

//MAC_3538 replaced by MAC_5827

//MAC_3537 replaced by MAC_5826

//MAC_3536 replaced by MAC_5827

//MAC_3535 replaced by MAC_5827

//MAC_3534 replaced by MAC_5826

//MAC_3545 replaced by MAC_5827

//MAC_3544 replaced by MAC_5827

//MAC_3543 replaced by MAC_5826

//MAC_3542 replaced by MAC_5827

//MAC_3541 replaced by MAC_5827

//MAC_3540 replaced by MAC_5826

//MAC_3551 replaced by MAC_5827

//MAC_3550 replaced by MAC_5827

//MAC_3549 replaced by MAC_5826

//MAC_3548 replaced by MAC_5827

//MAC_3547 replaced by MAC_5827

//MAC_3546 replaced by MAC_5826

//MAC_3557 replaced by MAC_5827

//MAC_3556 replaced by MAC_5827

//MAC_3555 replaced by MAC_5826

//MAC_3554 replaced by MAC_5827

//MAC_3553 replaced by MAC_5827

//MAC_3552 replaced by MAC_5826

//MAC_3563 replaced by MAC_5827

//MAC_3562 replaced by MAC_5827

//MAC_3561 replaced by MAC_5826

//MAC_3560 replaced by MAC_5827

//MAC_3559 replaced by MAC_5827

//MAC_3558 replaced by MAC_5826

//MAC_3569 replaced by MAC_5827

//MAC_3568 replaced by MAC_5827

//MAC_3567 replaced by MAC_5826

//MAC_3566 replaced by MAC_5827

//MAC_3565 replaced by MAC_5827

//MAC_3564 replaced by MAC_5826

//MAC_3575 replaced by MAC_5827

//MAC_3574 replaced by MAC_5827

//MAC_3573 replaced by MAC_5826

//MAC_3572 replaced by MAC_5827

//MAC_3571 replaced by MAC_5827

//MAC_3570 replaced by MAC_5826

//MAC_3581 replaced by MAC_5827

//MAC_3580 replaced by MAC_5827

//MAC_3579 replaced by MAC_5826

//MAC_3578 replaced by MAC_5827

//MAC_3577 replaced by MAC_5827

//MAC_3576 replaced by MAC_5826

//MAC_3587 replaced by MAC_5827

//MAC_3586 replaced by MAC_5827

//MAC_3585 replaced by MAC_5826

//MAC_3584 replaced by MAC_5827

//MAC_3583 replaced by MAC_5827

//MAC_3582 replaced by MAC_5826

//MAC_3593 replaced by MAC_5827

//MAC_3592 replaced by MAC_5827

//MAC_3591 replaced by MAC_5826

//MAC_3590 replaced by MAC_5827

//MAC_3589 replaced by MAC_5827

//MAC_3588 replaced by MAC_5826

//MAC_3599 replaced by MAC_5827

//MAC_3598 replaced by MAC_5827

//MAC_3597 replaced by MAC_5826

//MAC_3596 replaced by MAC_5827

//MAC_3595 replaced by MAC_5827

//MAC_3594 replaced by MAC_5826

//MAC_3605 replaced by MAC_5827

//MAC_3604 replaced by MAC_5827

//MAC_3603 replaced by MAC_5826

//MAC_3602 replaced by MAC_5827

//MAC_3601 replaced by MAC_5827

//MAC_3600 replaced by MAC_5826

//MAC_3611 replaced by MAC_5827

//MAC_3610 replaced by MAC_5827

//MAC_3609 replaced by MAC_5826

//MAC_3608 replaced by MAC_5827

//MAC_3607 replaced by MAC_5827

//MAC_3606 replaced by MAC_5826

//MAC_3617 replaced by MAC_5827

//MAC_3616 replaced by MAC_5827

//MAC_3615 replaced by MAC_5826

//MAC_3614 replaced by MAC_5827

//MAC_3613 replaced by MAC_5827

//MAC_3612 replaced by MAC_5826

//MAC_3623 replaced by MAC_5827

//MAC_3622 replaced by MAC_5827

//MAC_3621 replaced by MAC_5826

//MAC_3620 replaced by MAC_5827

//MAC_3619 replaced by MAC_5827

//MAC_3618 replaced by MAC_5826

//MAC_3629 replaced by MAC_5827

//MAC_3628 replaced by MAC_5827

//MAC_3627 replaced by MAC_5826

//MAC_3626 replaced by MAC_5827

//MAC_3625 replaced by MAC_5827

//MAC_3624 replaced by MAC_5826

//MAC_3635 replaced by MAC_5827

//MAC_3634 replaced by MAC_5827

//MAC_3633 replaced by MAC_5826

//MAC_3632 replaced by MAC_5827

//MAC_3631 replaced by MAC_5827

//MAC_3630 replaced by MAC_5826

//MAC_3641 replaced by MAC_5827

//MAC_3640 replaced by MAC_5827

//MAC_3639 replaced by MAC_5826

//MAC_3638 replaced by MAC_5827

//MAC_3637 replaced by MAC_5827

//MAC_3636 replaced by MAC_5826

//MAC_3647 replaced by MAC_5827

//MAC_3646 replaced by MAC_5827

//MAC_3645 replaced by MAC_5826

//MAC_3644 replaced by MAC_5827

//MAC_3643 replaced by MAC_5827

//MAC_3642 replaced by MAC_5826

//MAC_3653 replaced by MAC_5827

//MAC_3652 replaced by MAC_5827

//MAC_3651 replaced by MAC_5826

//MAC_3650 replaced by MAC_5827

//MAC_3649 replaced by MAC_5827

//MAC_3648 replaced by MAC_5826

//MAC_3659 replaced by MAC_5827

//MAC_3658 replaced by MAC_5827

//MAC_3657 replaced by MAC_5826

//MAC_3656 replaced by MAC_5827

//MAC_3655 replaced by MAC_5827

//MAC_3654 replaced by MAC_5826

//MAC_3665 replaced by MAC_5827

//MAC_3664 replaced by MAC_5827

//MAC_3663 replaced by MAC_5826

//MAC_3662 replaced by MAC_5827

//MAC_3661 replaced by MAC_5827

//MAC_3660 replaced by MAC_5826

//MAC_3671 replaced by MAC_5827

//MAC_3670 replaced by MAC_5827

//MAC_3669 replaced by MAC_5826

//MAC_3668 replaced by MAC_5827

//MAC_3667 replaced by MAC_5827

//MAC_3666 replaced by MAC_5826

//MAC_3677 replaced by MAC_5827

//MAC_3676 replaced by MAC_5827

//MAC_3675 replaced by MAC_5826

//MAC_3674 replaced by MAC_5827

//MAC_3673 replaced by MAC_5827

//MAC_3672 replaced by MAC_5826

//MAC_3683 replaced by MAC_5827

//MAC_3682 replaced by MAC_5827

//MAC_3681 replaced by MAC_5826

//MAC_3680 replaced by MAC_5827

//MAC_3679 replaced by MAC_5827

//MAC_3678 replaced by MAC_5826

//MAC_3689 replaced by MAC_5827

//MAC_3688 replaced by MAC_5827

//MAC_3687 replaced by MAC_5826

//MAC_3686 replaced by MAC_5827

//MAC_3685 replaced by MAC_5827

//MAC_3684 replaced by MAC_5826

//MAC_3695 replaced by MAC_5827

//MAC_3694 replaced by MAC_5827

//MAC_3693 replaced by MAC_5826

//MAC_3692 replaced by MAC_5827

//MAC_3691 replaced by MAC_5827

//MAC_3690 replaced by MAC_5826

//MAC_3701 replaced by MAC_5827

//MAC_3700 replaced by MAC_5827

//MAC_3699 replaced by MAC_5826

//MAC_3698 replaced by MAC_5827

//MAC_3697 replaced by MAC_5827

//MAC_3696 replaced by MAC_5826

//MAC_3707 replaced by MAC_5827

//MAC_3706 replaced by MAC_5827

//MAC_3705 replaced by MAC_5826

//MAC_3704 replaced by MAC_5827

//MAC_3703 replaced by MAC_5827

//MAC_3702 replaced by MAC_5826

//MAC_3713 replaced by MAC_5827

//MAC_3712 replaced by MAC_5827

//MAC_3711 replaced by MAC_5826

//MAC_3710 replaced by MAC_5827

//MAC_3709 replaced by MAC_5827

//MAC_3708 replaced by MAC_5826

//MAC_3719 replaced by MAC_5827

//MAC_3718 replaced by MAC_5827

//MAC_3717 replaced by MAC_5826

//MAC_3716 replaced by MAC_5827

//MAC_3715 replaced by MAC_5827

//MAC_3714 replaced by MAC_5826

//MAC_3725 replaced by MAC_5827

//MAC_3724 replaced by MAC_5827

//MAC_3723 replaced by MAC_5826

//MAC_3722 replaced by MAC_5827

//MAC_3721 replaced by MAC_5827

//MAC_3720 replaced by MAC_5826

//MAC_3731 replaced by MAC_5827

//MAC_3730 replaced by MAC_5827

//MAC_3729 replaced by MAC_5826

//MAC_3728 replaced by MAC_5827

//MAC_3727 replaced by MAC_5827

//MAC_3726 replaced by MAC_5826

//MAC_3737 replaced by MAC_5827

//MAC_3736 replaced by MAC_5827

//MAC_3735 replaced by MAC_5826

//MAC_3734 replaced by MAC_5827

//MAC_3733 replaced by MAC_5827

//MAC_3732 replaced by MAC_5826

//MAC_3743 replaced by MAC_5827

//MAC_3742 replaced by MAC_5827

//MAC_3741 replaced by MAC_5826

//MAC_3740 replaced by MAC_5827

//MAC_3739 replaced by MAC_5827

//MAC_3738 replaced by MAC_5826

//MAC_3749 replaced by MAC_5827

//MAC_3748 replaced by MAC_5827

//MAC_3747 replaced by MAC_5826

//MAC_3746 replaced by MAC_5827

//MAC_3745 replaced by MAC_5827

//MAC_3744 replaced by MAC_5826

//MAC_3755 replaced by MAC_5827

//MAC_3754 replaced by MAC_5827

//MAC_3753 replaced by MAC_5826

//MAC_3752 replaced by MAC_5827

//MAC_3751 replaced by MAC_5827

//MAC_3750 replaced by MAC_5826

//MAC_3761 replaced by MAC_5827

//MAC_3760 replaced by MAC_5827

//MAC_3759 replaced by MAC_5826

//MAC_3758 replaced by MAC_5827

//MAC_3757 replaced by MAC_5827

//MAC_3756 replaced by MAC_5826

//MAC_3767 replaced by MAC_5827

//MAC_3766 replaced by MAC_5827

//MAC_3765 replaced by MAC_5826

//MAC_3764 replaced by MAC_5827

//MAC_3763 replaced by MAC_5827

//MAC_3762 replaced by MAC_5826

//MAC_3773 replaced by MAC_5827

//MAC_3772 replaced by MAC_5827

//MAC_3771 replaced by MAC_5826

//MAC_3770 replaced by MAC_5827

//MAC_3769 replaced by MAC_5827

//MAC_3768 replaced by MAC_5826

//MAC_3779 replaced by MAC_5827

//MAC_3778 replaced by MAC_5827

//MAC_3777 replaced by MAC_5826

//MAC_3776 replaced by MAC_5827

//MAC_3775 replaced by MAC_5827

//MAC_3774 replaced by MAC_5826

//MAC_3785 replaced by MAC_5827

//MAC_3784 replaced by MAC_5827

//MAC_3783 replaced by MAC_5826

//MAC_3782 replaced by MAC_5827

//MAC_3781 replaced by MAC_5827

//MAC_3780 replaced by MAC_5826

//MAC_3791 replaced by MAC_5827

//MAC_3790 replaced by MAC_5827

//MAC_3789 replaced by MAC_5826

//MAC_3788 replaced by MAC_5827

//MAC_3787 replaced by MAC_5827

//MAC_3786 replaced by MAC_5826

//MAC_3797 replaced by MAC_5827

//MAC_3796 replaced by MAC_5827

//MAC_3795 replaced by MAC_5826

//MAC_3794 replaced by MAC_5827

//MAC_3793 replaced by MAC_5827

//MAC_3792 replaced by MAC_5826

//MAC_3803 replaced by MAC_5827

//MAC_3802 replaced by MAC_5827

//MAC_3801 replaced by MAC_5826

//MAC_3800 replaced by MAC_5827

//MAC_3799 replaced by MAC_5827

//MAC_3798 replaced by MAC_5826

//MAC_3809 replaced by MAC_5827

//MAC_3808 replaced by MAC_5827

//MAC_3807 replaced by MAC_5826

//MAC_3806 replaced by MAC_5827

//MAC_3805 replaced by MAC_5827

//MAC_3804 replaced by MAC_5826

//MAC_3815 replaced by MAC_5827

//MAC_3814 replaced by MAC_5827

//MAC_3813 replaced by MAC_5826

//MAC_3812 replaced by MAC_5827

//MAC_3811 replaced by MAC_5827

//MAC_3810 replaced by MAC_5826

//MAC_3821 replaced by MAC_5827

//MAC_3820 replaced by MAC_5827

//MAC_3819 replaced by MAC_5826

//MAC_3818 replaced by MAC_5827

//MAC_3817 replaced by MAC_5827

//MAC_3816 replaced by MAC_5826

//MAC_3827 replaced by MAC_5827

//MAC_3826 replaced by MAC_5827

//MAC_3825 replaced by MAC_5826

//MAC_3824 replaced by MAC_5827

//MAC_3823 replaced by MAC_5827

//MAC_3822 replaced by MAC_5826

//MAC_3833 replaced by MAC_5827

//MAC_3832 replaced by MAC_5827

//MAC_3831 replaced by MAC_5826

//MAC_3830 replaced by MAC_5827

//MAC_3829 replaced by MAC_5827

//MAC_3828 replaced by MAC_5826

//MAC_3839 replaced by MAC_5827

//MAC_3838 replaced by MAC_5827

//MAC_3837 replaced by MAC_5826

//MAC_3836 replaced by MAC_5827

//MAC_3835 replaced by MAC_5827

//MAC_3834 replaced by MAC_5826

//MAC_3845 replaced by MAC_5827

//MAC_3844 replaced by MAC_5827

//MAC_3843 replaced by MAC_5826

//MAC_3842 replaced by MAC_5827

//MAC_3841 replaced by MAC_5827

//MAC_3840 replaced by MAC_5826

//MAC_3851 replaced by MAC_5827

//MAC_3850 replaced by MAC_5827

//MAC_3849 replaced by MAC_5826

//MAC_3848 replaced by MAC_5827

//MAC_3847 replaced by MAC_5827

//MAC_3846 replaced by MAC_5826

//MAC_3857 replaced by MAC_5827

//MAC_3856 replaced by MAC_5827

//MAC_3855 replaced by MAC_5826

//MAC_3854 replaced by MAC_5827

//MAC_3853 replaced by MAC_5827

//MAC_3852 replaced by MAC_5826

//MAC_3863 replaced by MAC_5827

//MAC_3862 replaced by MAC_5827

//MAC_3861 replaced by MAC_5826

//MAC_3860 replaced by MAC_5827

//MAC_3859 replaced by MAC_5827

//MAC_3858 replaced by MAC_5826

//MAC_3869 replaced by MAC_5827

//MAC_3868 replaced by MAC_5827

//MAC_3867 replaced by MAC_5826

//MAC_3866 replaced by MAC_5827

//MAC_3865 replaced by MAC_5827

//MAC_3864 replaced by MAC_5826

//MAC_3875 replaced by MAC_5827

//MAC_3874 replaced by MAC_5827

//MAC_3873 replaced by MAC_5826

//MAC_3872 replaced by MAC_5827

//MAC_3871 replaced by MAC_5827

//MAC_3870 replaced by MAC_5826

//MAC_3881 replaced by MAC_5827

//MAC_3880 replaced by MAC_5827

//MAC_3879 replaced by MAC_5826

//MAC_3878 replaced by MAC_5827

//MAC_3877 replaced by MAC_5827

//MAC_3876 replaced by MAC_5826

//MAC_3887 replaced by MAC_5827

//MAC_3886 replaced by MAC_5827

//MAC_3885 replaced by MAC_5826

//MAC_3884 replaced by MAC_5827

//MAC_3883 replaced by MAC_5827

//MAC_3882 replaced by MAC_5826

//MAC_3893 replaced by MAC_5827

//MAC_3892 replaced by MAC_5827

//MAC_3891 replaced by MAC_5826

//MAC_3890 replaced by MAC_5827

//MAC_3889 replaced by MAC_5827

//MAC_3888 replaced by MAC_5826

//MAC_3899 replaced by MAC_5827

//MAC_3898 replaced by MAC_5827

//MAC_3897 replaced by MAC_5826

//MAC_3896 replaced by MAC_5827

//MAC_3895 replaced by MAC_5827

//MAC_3894 replaced by MAC_5826

//MAC_3905 replaced by MAC_5827

//MAC_3904 replaced by MAC_5827

//MAC_3903 replaced by MAC_5826

//MAC_3902 replaced by MAC_5827

//MAC_3901 replaced by MAC_5827

//MAC_3900 replaced by MAC_5826

//MAC_3911 replaced by MAC_5827

//MAC_3910 replaced by MAC_5827

//MAC_3909 replaced by MAC_5826

//MAC_3908 replaced by MAC_5827

//MAC_3907 replaced by MAC_5827

//MAC_3906 replaced by MAC_5826

//MAC_3917 replaced by MAC_5827

//MAC_3916 replaced by MAC_5827

//MAC_3915 replaced by MAC_5826

//MAC_3914 replaced by MAC_5827

//MAC_3913 replaced by MAC_5827

//MAC_3912 replaced by MAC_5826

//MAC_3923 replaced by MAC_5827

//MAC_3922 replaced by MAC_5827

//MAC_3921 replaced by MAC_5826

//MAC_3920 replaced by MAC_5827

//MAC_3919 replaced by MAC_5827

//MAC_3918 replaced by MAC_5826

//MAC_3929 replaced by MAC_5827

//MAC_3928 replaced by MAC_5827

//MAC_3927 replaced by MAC_5826

//MAC_3926 replaced by MAC_5827

//MAC_3925 replaced by MAC_5827

//MAC_3924 replaced by MAC_5826

//MAC_3935 replaced by MAC_5827

//MAC_3934 replaced by MAC_5827

//MAC_3933 replaced by MAC_5826

//MAC_3932 replaced by MAC_5827

//MAC_3931 replaced by MAC_5827

//MAC_3930 replaced by MAC_5826

//MAC_3941 replaced by MAC_5827

//MAC_3940 replaced by MAC_5827

//MAC_3939 replaced by MAC_5826

//MAC_3938 replaced by MAC_5827

//MAC_3937 replaced by MAC_5827

//MAC_3936 replaced by MAC_5826

//MAC_3947 replaced by MAC_5827

//MAC_3946 replaced by MAC_5827

//MAC_3945 replaced by MAC_5826

//MAC_3944 replaced by MAC_5827

//MAC_3943 replaced by MAC_5827

//MAC_3942 replaced by MAC_5826

//MAC_3953 replaced by MAC_5827

//MAC_3952 replaced by MAC_5827

//MAC_3951 replaced by MAC_5826

//MAC_3950 replaced by MAC_5827

//MAC_3949 replaced by MAC_5827

//MAC_3948 replaced by MAC_5826

//MAC_3959 replaced by MAC_5827

//MAC_3958 replaced by MAC_5827

//MAC_3957 replaced by MAC_5826

//MAC_3956 replaced by MAC_5827

//MAC_3955 replaced by MAC_5827

//MAC_3954 replaced by MAC_5826

//MAC_3965 replaced by MAC_5827

//MAC_3964 replaced by MAC_5827

//MAC_3963 replaced by MAC_5826

//MAC_3962 replaced by MAC_5827

//MAC_3961 replaced by MAC_5827

//MAC_3960 replaced by MAC_5826

//MAC_3971 replaced by MAC_5827

//MAC_3970 replaced by MAC_5827

//MAC_3969 replaced by MAC_5826

//MAC_3968 replaced by MAC_5827

//MAC_3967 replaced by MAC_5827

//MAC_3966 replaced by MAC_5826

//MAC_3977 replaced by MAC_5827

//MAC_3976 replaced by MAC_5827

//MAC_3975 replaced by MAC_5826

//MAC_3974 replaced by MAC_5827

//MAC_3973 replaced by MAC_5827

//MAC_3972 replaced by MAC_5826

//MAC_3983 replaced by MAC_5827

//MAC_3982 replaced by MAC_5827

//MAC_3981 replaced by MAC_5826

//MAC_3980 replaced by MAC_5827

//MAC_3979 replaced by MAC_5827

//MAC_3978 replaced by MAC_5826

//MAC_3989 replaced by MAC_5827

//MAC_3988 replaced by MAC_5827

//MAC_3987 replaced by MAC_5826

//MAC_3986 replaced by MAC_5827

//MAC_3985 replaced by MAC_5827

//MAC_3984 replaced by MAC_5826

//MAC_3995 replaced by MAC_5827

//MAC_3994 replaced by MAC_5827

//MAC_3993 replaced by MAC_5826

//MAC_3992 replaced by MAC_5827

//MAC_3991 replaced by MAC_5827

//MAC_3990 replaced by MAC_5826

//MAC_4001 replaced by MAC_5827

//MAC_4000 replaced by MAC_5827

//MAC_3999 replaced by MAC_5826

//MAC_3998 replaced by MAC_5827

//MAC_3997 replaced by MAC_5827

//MAC_3996 replaced by MAC_5826

//MAC_4007 replaced by MAC_5827

//MAC_4006 replaced by MAC_5827

//MAC_4005 replaced by MAC_5826

//MAC_4004 replaced by MAC_5827

//MAC_4003 replaced by MAC_5827

//MAC_4002 replaced by MAC_5826

//MAC_4013 replaced by MAC_5827

//MAC_4012 replaced by MAC_5827

//MAC_4011 replaced by MAC_5826

//MAC_4010 replaced by MAC_5827

//MAC_4009 replaced by MAC_5827

//MAC_4008 replaced by MAC_5826

//MAC_4019 replaced by MAC_5827

//MAC_4018 replaced by MAC_5827

//MAC_4017 replaced by MAC_5826

//MAC_4016 replaced by MAC_5827

//MAC_4015 replaced by MAC_5827

//MAC_4014 replaced by MAC_5826

//MAC_4025 replaced by MAC_5827

//MAC_4024 replaced by MAC_5827

//MAC_4023 replaced by MAC_5826

//MAC_4022 replaced by MAC_5827

//MAC_4021 replaced by MAC_5827

//MAC_4020 replaced by MAC_5826

//MAC_4031 replaced by MAC_5827

//MAC_4030 replaced by MAC_5827

//MAC_4029 replaced by MAC_5826

//MAC_4028 replaced by MAC_5827

//MAC_4027 replaced by MAC_5827

//MAC_4026 replaced by MAC_5826

//MAC_4037 replaced by MAC_5827

//MAC_4036 replaced by MAC_5827

//MAC_4035 replaced by MAC_5826

//MAC_4034 replaced by MAC_5827

//MAC_4033 replaced by MAC_5827

//MAC_4032 replaced by MAC_5826

//MAC_4043 replaced by MAC_5827

//MAC_4042 replaced by MAC_5827

//MAC_4041 replaced by MAC_5826

//MAC_4040 replaced by MAC_5827

//MAC_4039 replaced by MAC_5827

//MAC_4038 replaced by MAC_5826

//MAC_4049 replaced by MAC_5827

//MAC_4048 replaced by MAC_5827

//MAC_4047 replaced by MAC_5826

//MAC_4046 replaced by MAC_5827

//MAC_4045 replaced by MAC_5827

//MAC_4044 replaced by MAC_5826

//MAC_4055 replaced by MAC_5827

//MAC_4054 replaced by MAC_5827

//MAC_4053 replaced by MAC_5826

//MAC_4052 replaced by MAC_5827

//MAC_4051 replaced by MAC_5827

//MAC_4050 replaced by MAC_5826

//MAC_4061 replaced by MAC_5827

//MAC_4060 replaced by MAC_5827

//MAC_4059 replaced by MAC_5826

//MAC_4058 replaced by MAC_5827

//MAC_4057 replaced by MAC_5827

//MAC_4056 replaced by MAC_5826

//MAC_4067 replaced by MAC_5827

//MAC_4066 replaced by MAC_5827

//MAC_4065 replaced by MAC_5826

//MAC_4064 replaced by MAC_5827

//MAC_4063 replaced by MAC_5827

//MAC_4062 replaced by MAC_5826

//MAC_4073 replaced by MAC_5827

//MAC_4072 replaced by MAC_5827

//MAC_4071 replaced by MAC_5826

//MAC_4070 replaced by MAC_5827

//MAC_4069 replaced by MAC_5827

//MAC_4068 replaced by MAC_5826

//MAC_4079 replaced by MAC_5827

//MAC_4078 replaced by MAC_5827

//MAC_4077 replaced by MAC_5826

//MAC_4076 replaced by MAC_5827

//MAC_4075 replaced by MAC_5827

//MAC_4074 replaced by MAC_5826

//MAC_4085 replaced by MAC_5827

//MAC_4084 replaced by MAC_5827

//MAC_4083 replaced by MAC_5826

//MAC_4082 replaced by MAC_5827

//MAC_4081 replaced by MAC_5827

//MAC_4080 replaced by MAC_5826

//MAC_4091 replaced by MAC_5827

//MAC_4090 replaced by MAC_5827

//MAC_4089 replaced by MAC_5826

//MAC_4088 replaced by MAC_5827

//MAC_4087 replaced by MAC_5827

//MAC_4086 replaced by MAC_5826

//MAC_4097 replaced by MAC_5827

//MAC_4096 replaced by MAC_5827

//MAC_4095 replaced by MAC_5826

//MAC_4094 replaced by MAC_5827

//MAC_4093 replaced by MAC_5827

//MAC_4092 replaced by MAC_5826

//MAC_4103 replaced by MAC_5827

//MAC_4102 replaced by MAC_5827

//MAC_4101 replaced by MAC_5826

//MAC_4100 replaced by MAC_5827

//MAC_4099 replaced by MAC_5827

//MAC_4098 replaced by MAC_5826

//MAC_4109 replaced by MAC_5827

//MAC_4108 replaced by MAC_5827

//MAC_4107 replaced by MAC_5826

//MAC_4106 replaced by MAC_5827

//MAC_4105 replaced by MAC_5827

//MAC_4104 replaced by MAC_5826

//MAC_4115 replaced by MAC_5827

//MAC_4114 replaced by MAC_5827

//MAC_4113 replaced by MAC_5826

//MAC_4112 replaced by MAC_5827

//MAC_4111 replaced by MAC_5827

//MAC_4110 replaced by MAC_5826

//MAC_4121 replaced by MAC_5827

//MAC_4120 replaced by MAC_5827

//MAC_4119 replaced by MAC_5826

//MAC_4118 replaced by MAC_5827

//MAC_4117 replaced by MAC_5827

//MAC_4116 replaced by MAC_5826

//MAC_4127 replaced by MAC_5827

//MAC_4126 replaced by MAC_5827

//MAC_4125 replaced by MAC_5826

//MAC_4124 replaced by MAC_5827

//MAC_4123 replaced by MAC_5827

//MAC_4122 replaced by MAC_5826

//MAC_4133 replaced by MAC_5827

//MAC_4132 replaced by MAC_5827

//MAC_4131 replaced by MAC_5826

//MAC_4130 replaced by MAC_5827

//MAC_4129 replaced by MAC_5827

//MAC_4128 replaced by MAC_5826

//MAC_4139 replaced by MAC_5827

//MAC_4138 replaced by MAC_5827

//MAC_4137 replaced by MAC_5826

//MAC_4136 replaced by MAC_5827

//MAC_4135 replaced by MAC_5827

//MAC_4134 replaced by MAC_5826

//MAC_4145 replaced by MAC_5827

//MAC_4144 replaced by MAC_5827

//MAC_4143 replaced by MAC_5826

//MAC_4142 replaced by MAC_5827

//MAC_4141 replaced by MAC_5827

//MAC_4140 replaced by MAC_5826

//MAC_4151 replaced by MAC_5827

//MAC_4150 replaced by MAC_5827

//MAC_4149 replaced by MAC_5826

//MAC_4148 replaced by MAC_5827

//MAC_4147 replaced by MAC_5827

//MAC_4146 replaced by MAC_5826

//MAC_4157 replaced by MAC_5827

//MAC_4156 replaced by MAC_5827

//MAC_4155 replaced by MAC_5826

//MAC_4154 replaced by MAC_5827

//MAC_4153 replaced by MAC_5827

//MAC_4152 replaced by MAC_5826

//MAC_4163 replaced by MAC_5827

//MAC_4162 replaced by MAC_5827

//MAC_4161 replaced by MAC_5826

//MAC_4160 replaced by MAC_5827

//MAC_4159 replaced by MAC_5827

//MAC_4158 replaced by MAC_5826

//MAC_4169 replaced by MAC_5827

//MAC_4168 replaced by MAC_5827

//MAC_4167 replaced by MAC_5826

//MAC_4166 replaced by MAC_5827

//MAC_4165 replaced by MAC_5827

//MAC_4164 replaced by MAC_5826

//MAC_4175 replaced by MAC_5827

//MAC_4174 replaced by MAC_5827

//MAC_4173 replaced by MAC_5826

//MAC_4172 replaced by MAC_5827

//MAC_4171 replaced by MAC_5827

//MAC_4170 replaced by MAC_5826

//MAC_4181 replaced by MAC_5827

//MAC_4180 replaced by MAC_5827

//MAC_4179 replaced by MAC_5826

//MAC_4178 replaced by MAC_5827

//MAC_4177 replaced by MAC_5827

//MAC_4176 replaced by MAC_5826

//MAC_4187 replaced by MAC_5827

//MAC_4186 replaced by MAC_5827

//MAC_4185 replaced by MAC_5826

//MAC_4184 replaced by MAC_5827

//MAC_4183 replaced by MAC_5827

//MAC_4182 replaced by MAC_5826

//MAC_4193 replaced by MAC_5827

//MAC_4192 replaced by MAC_5827

//MAC_4191 replaced by MAC_5826

//MAC_4190 replaced by MAC_5827

//MAC_4189 replaced by MAC_5827

//MAC_4188 replaced by MAC_5826

//MAC_4199 replaced by MAC_5827

//MAC_4198 replaced by MAC_5827

//MAC_4197 replaced by MAC_5826

//MAC_4196 replaced by MAC_5827

//MAC_4195 replaced by MAC_5827

//MAC_4194 replaced by MAC_5826

//MAC_4205 replaced by MAC_5827

//MAC_4204 replaced by MAC_5827

//MAC_4203 replaced by MAC_5826

//MAC_4202 replaced by MAC_5827

//MAC_4201 replaced by MAC_5827

//MAC_4200 replaced by MAC_5826

//MAC_4211 replaced by MAC_5827

//MAC_4210 replaced by MAC_5827

//MAC_4209 replaced by MAC_5826

//MAC_4208 replaced by MAC_5827

//MAC_4207 replaced by MAC_5827

//MAC_4206 replaced by MAC_5826

//MAC_4217 replaced by MAC_5827

//MAC_4216 replaced by MAC_5827

//MAC_4215 replaced by MAC_5826

//MAC_4214 replaced by MAC_5827

//MAC_4213 replaced by MAC_5827

//MAC_4212 replaced by MAC_5826

//MAC_4223 replaced by MAC_5827

//MAC_4222 replaced by MAC_5827

//MAC_4221 replaced by MAC_5826

//MAC_4220 replaced by MAC_5827

//MAC_4219 replaced by MAC_5827

//MAC_4218 replaced by MAC_5826

//MAC_4229 replaced by MAC_5827

//MAC_4228 replaced by MAC_5827

//MAC_4227 replaced by MAC_5826

//MAC_4226 replaced by MAC_5827

//MAC_4225 replaced by MAC_5827

//MAC_4224 replaced by MAC_5826

//MAC_4235 replaced by MAC_5827

//MAC_4234 replaced by MAC_5827

//MAC_4233 replaced by MAC_5826

//MAC_4232 replaced by MAC_5827

//MAC_4231 replaced by MAC_5827

//MAC_4230 replaced by MAC_5826

//MAC_4241 replaced by MAC_5827

//MAC_4240 replaced by MAC_5827

//MAC_4239 replaced by MAC_5826

//MAC_4238 replaced by MAC_5827

//MAC_4237 replaced by MAC_5827

//MAC_4236 replaced by MAC_5826

//MAC_4247 replaced by MAC_5827

//MAC_4246 replaced by MAC_5827

//MAC_4245 replaced by MAC_5826

//MAC_4244 replaced by MAC_5827

//MAC_4243 replaced by MAC_5827

//MAC_4242 replaced by MAC_5826

//MAC_4253 replaced by MAC_5827

//MAC_4252 replaced by MAC_5827

//MAC_4251 replaced by MAC_5826

//MAC_4250 replaced by MAC_5827

//MAC_4249 replaced by MAC_5827

//MAC_4248 replaced by MAC_5826

//MAC_4259 replaced by MAC_5827

//MAC_4258 replaced by MAC_5827

//MAC_4257 replaced by MAC_5826

//MAC_4256 replaced by MAC_5827

//MAC_4255 replaced by MAC_5827

//MAC_4254 replaced by MAC_5826

//MAC_4265 replaced by MAC_5827

//MAC_4264 replaced by MAC_5827

//MAC_4263 replaced by MAC_5826

//MAC_4262 replaced by MAC_5827

//MAC_4261 replaced by MAC_5827

//MAC_4260 replaced by MAC_5826

//MAC_4271 replaced by MAC_5827

//MAC_4270 replaced by MAC_5827

//MAC_4269 replaced by MAC_5826

//MAC_4268 replaced by MAC_5827

//MAC_4267 replaced by MAC_5827

//MAC_4266 replaced by MAC_5826

//MAC_4277 replaced by MAC_5827

//MAC_4276 replaced by MAC_5827

//MAC_4275 replaced by MAC_5826

//MAC_4274 replaced by MAC_5827

//MAC_4273 replaced by MAC_5827

//MAC_4272 replaced by MAC_5826

//MAC_4283 replaced by MAC_5827

//MAC_4282 replaced by MAC_5827

//MAC_4281 replaced by MAC_5826

//MAC_4280 replaced by MAC_5827

//MAC_4279 replaced by MAC_5827

//MAC_4278 replaced by MAC_5826

//MAC_4289 replaced by MAC_5827

//MAC_4288 replaced by MAC_5827

//MAC_4287 replaced by MAC_5826

//MAC_4286 replaced by MAC_5827

//MAC_4285 replaced by MAC_5827

//MAC_4284 replaced by MAC_5826

//MAC_4295 replaced by MAC_5827

//MAC_4294 replaced by MAC_5827

//MAC_4293 replaced by MAC_5826

//MAC_4292 replaced by MAC_5827

//MAC_4291 replaced by MAC_5827

//MAC_4290 replaced by MAC_5826

//MAC_4301 replaced by MAC_5827

//MAC_4300 replaced by MAC_5827

//MAC_4299 replaced by MAC_5826

//MAC_4298 replaced by MAC_5827

//MAC_4297 replaced by MAC_5827

//MAC_4296 replaced by MAC_5826

//MAC_4307 replaced by MAC_5827

//MAC_4306 replaced by MAC_5827

//MAC_4305 replaced by MAC_5826

//MAC_4304 replaced by MAC_5827

//MAC_4303 replaced by MAC_5827

//MAC_4302 replaced by MAC_5826

//MAC_4313 replaced by MAC_5827

//MAC_4312 replaced by MAC_5827

//MAC_4311 replaced by MAC_5826

//MAC_4310 replaced by MAC_5827

//MAC_4309 replaced by MAC_5827

//MAC_4308 replaced by MAC_5826

//MAC_4319 replaced by MAC_5827

//MAC_4318 replaced by MAC_5827

//MAC_4317 replaced by MAC_5826

//MAC_4316 replaced by MAC_5827

//MAC_4315 replaced by MAC_5827

//MAC_4314 replaced by MAC_5826

//MAC_4325 replaced by MAC_5827

//MAC_4324 replaced by MAC_5827

//MAC_4323 replaced by MAC_5826

//MAC_4322 replaced by MAC_5827

//MAC_4321 replaced by MAC_5827

//MAC_4320 replaced by MAC_5826

//MAC_4331 replaced by MAC_5827

//MAC_4330 replaced by MAC_5827

//MAC_4329 replaced by MAC_5826

//MAC_4328 replaced by MAC_5827

//MAC_4327 replaced by MAC_5827

//MAC_4326 replaced by MAC_5826

//MAC_4337 replaced by MAC_5827

//MAC_4336 replaced by MAC_5827

//MAC_4335 replaced by MAC_5826

//MAC_4334 replaced by MAC_5827

//MAC_4333 replaced by MAC_5827

//MAC_4332 replaced by MAC_5826

//MAC_4343 replaced by MAC_5827

//MAC_4342 replaced by MAC_5827

//MAC_4341 replaced by MAC_5826

//MAC_4340 replaced by MAC_5827

//MAC_4339 replaced by MAC_5827

//MAC_4338 replaced by MAC_5826

//MAC_4349 replaced by MAC_5827

//MAC_4348 replaced by MAC_5827

//MAC_4347 replaced by MAC_5826

//MAC_4346 replaced by MAC_5827

//MAC_4345 replaced by MAC_5827

//MAC_4344 replaced by MAC_5826

//MAC_4355 replaced by MAC_5827

//MAC_4354 replaced by MAC_5827

//MAC_4353 replaced by MAC_5826

//MAC_4352 replaced by MAC_5827

//MAC_4351 replaced by MAC_5827

//MAC_4350 replaced by MAC_5826

//MAC_4361 replaced by MAC_5827

//MAC_4360 replaced by MAC_5827

//MAC_4359 replaced by MAC_5826

//MAC_4358 replaced by MAC_5827

//MAC_4357 replaced by MAC_5827

//MAC_4356 replaced by MAC_5826

//MAC_4367 replaced by MAC_5827

//MAC_4366 replaced by MAC_5827

//MAC_4365 replaced by MAC_5826

//MAC_4364 replaced by MAC_5827

//MAC_4363 replaced by MAC_5827

//MAC_4362 replaced by MAC_5826

//MAC_4373 replaced by MAC_5827

//MAC_4372 replaced by MAC_5827

//MAC_4371 replaced by MAC_5826

//MAC_4370 replaced by MAC_5827

//MAC_4369 replaced by MAC_5827

//MAC_4368 replaced by MAC_5826

//MAC_4379 replaced by MAC_5827

//MAC_4378 replaced by MAC_5827

//MAC_4377 replaced by MAC_5826

//MAC_4376 replaced by MAC_5827

//MAC_4375 replaced by MAC_5827

//MAC_4374 replaced by MAC_5826

//MAC_4385 replaced by MAC_5827

//MAC_4384 replaced by MAC_5827

//MAC_4383 replaced by MAC_5826

//MAC_4382 replaced by MAC_5827

//MAC_4381 replaced by MAC_5827

//MAC_4380 replaced by MAC_5826

//MAC_4391 replaced by MAC_5827

//MAC_4390 replaced by MAC_5827

//MAC_4389 replaced by MAC_5826

//MAC_4388 replaced by MAC_5827

//MAC_4387 replaced by MAC_5827

//MAC_4386 replaced by MAC_5826

//MAC_4397 replaced by MAC_5827

//MAC_4396 replaced by MAC_5827

//MAC_4395 replaced by MAC_5826

//MAC_4394 replaced by MAC_5827

//MAC_4393 replaced by MAC_5827

//MAC_4392 replaced by MAC_5826

//MAC_4403 replaced by MAC_5827

//MAC_4402 replaced by MAC_5827

//MAC_4401 replaced by MAC_5826

//MAC_4400 replaced by MAC_5827

//MAC_4399 replaced by MAC_5827

//MAC_4398 replaced by MAC_5826

//MAC_4409 replaced by MAC_5827

//MAC_4408 replaced by MAC_5827

//MAC_4407 replaced by MAC_5826

//MAC_4406 replaced by MAC_5827

//MAC_4405 replaced by MAC_5827

//MAC_4404 replaced by MAC_5826

//MAC_4415 replaced by MAC_5827

//MAC_4414 replaced by MAC_5827

//MAC_4413 replaced by MAC_5826

//MAC_4412 replaced by MAC_5827

//MAC_4411 replaced by MAC_5827

//MAC_4410 replaced by MAC_5826

//MAC_4421 replaced by MAC_5827

//MAC_4420 replaced by MAC_5827

//MAC_4419 replaced by MAC_5826

//MAC_4418 replaced by MAC_5827

//MAC_4417 replaced by MAC_5827

//MAC_4416 replaced by MAC_5826

//MAC_4427 replaced by MAC_5827

//MAC_4426 replaced by MAC_5827

//MAC_4425 replaced by MAC_5826

//MAC_4424 replaced by MAC_5827

//MAC_4423 replaced by MAC_5827

//MAC_4422 replaced by MAC_5826

//MAC_4433 replaced by MAC_5827

//MAC_4432 replaced by MAC_5827

//MAC_4431 replaced by MAC_5826

//MAC_4430 replaced by MAC_5827

//MAC_4429 replaced by MAC_5827

//MAC_4428 replaced by MAC_5826

//MAC_4439 replaced by MAC_5827

//MAC_4438 replaced by MAC_5827

//MAC_4437 replaced by MAC_5826

//MAC_4436 replaced by MAC_5827

//MAC_4435 replaced by MAC_5827

//MAC_4434 replaced by MAC_5826

//MAC_4445 replaced by MAC_5827

//MAC_4444 replaced by MAC_5827

//MAC_4443 replaced by MAC_5826

//MAC_4442 replaced by MAC_5827

//MAC_4441 replaced by MAC_5827

//MAC_4440 replaced by MAC_5826

//MAC_4451 replaced by MAC_5827

//MAC_4450 replaced by MAC_5827

//MAC_4449 replaced by MAC_5826

//MAC_4448 replaced by MAC_5827

//MAC_4447 replaced by MAC_5827

//MAC_4446 replaced by MAC_5826

//MAC_4457 replaced by MAC_5827

//MAC_4456 replaced by MAC_5827

//MAC_4455 replaced by MAC_5826

//MAC_4454 replaced by MAC_5827

//MAC_4453 replaced by MAC_5827

//MAC_4452 replaced by MAC_5826

//MAC_4463 replaced by MAC_5827

//MAC_4462 replaced by MAC_5827

//MAC_4461 replaced by MAC_5826

//MAC_4460 replaced by MAC_5827

//MAC_4459 replaced by MAC_5827

//MAC_4458 replaced by MAC_5826

//MAC_4469 replaced by MAC_5827

//MAC_4468 replaced by MAC_5827

//MAC_4467 replaced by MAC_5826

//MAC_4466 replaced by MAC_5827

//MAC_4465 replaced by MAC_5827

//MAC_4464 replaced by MAC_5826

//MAC_4475 replaced by MAC_5827

//MAC_4474 replaced by MAC_5827

//MAC_4473 replaced by MAC_5826

//MAC_4472 replaced by MAC_5827

//MAC_4471 replaced by MAC_5827

//MAC_4470 replaced by MAC_5826

//MAC_4481 replaced by MAC_5827

//MAC_4480 replaced by MAC_5827

//MAC_4479 replaced by MAC_5826

//MAC_4478 replaced by MAC_5827

//MAC_4477 replaced by MAC_5827

//MAC_4476 replaced by MAC_5826

//MAC_4487 replaced by MAC_5827

//MAC_4486 replaced by MAC_5827

//MAC_4485 replaced by MAC_5826

//MAC_4484 replaced by MAC_5827

//MAC_4483 replaced by MAC_5827

//MAC_4482 replaced by MAC_5826

//MAC_4493 replaced by MAC_5827

//MAC_4492 replaced by MAC_5827

//MAC_4491 replaced by MAC_5826

//MAC_4490 replaced by MAC_5827

//MAC_4489 replaced by MAC_5827

//MAC_4488 replaced by MAC_5826

//MAC_4499 replaced by MAC_5827

//MAC_4498 replaced by MAC_5827

//MAC_4497 replaced by MAC_5826

//MAC_4496 replaced by MAC_5827

//MAC_4495 replaced by MAC_5827

//MAC_4494 replaced by MAC_5826

//MAC_4505 replaced by MAC_5827

//MAC_4504 replaced by MAC_5827

//MAC_4503 replaced by MAC_5826

//MAC_4502 replaced by MAC_5827

//MAC_4501 replaced by MAC_5827

//MAC_4500 replaced by MAC_5826

//MAC_4511 replaced by MAC_5827

//MAC_4510 replaced by MAC_5827

//MAC_4509 replaced by MAC_5826

//MAC_4508 replaced by MAC_5827

//MAC_4507 replaced by MAC_5827

//MAC_4506 replaced by MAC_5826

//MAC_4517 replaced by MAC_5827

//MAC_4516 replaced by MAC_5827

//MAC_4515 replaced by MAC_5826

//MAC_4514 replaced by MAC_5827

//MAC_4513 replaced by MAC_5827

//MAC_4512 replaced by MAC_5826

//MAC_4523 replaced by MAC_5827

//MAC_4522 replaced by MAC_5827

//MAC_4521 replaced by MAC_5826

//MAC_4520 replaced by MAC_5827

//MAC_4519 replaced by MAC_5827

//MAC_4518 replaced by MAC_5826

//MAC_4529 replaced by MAC_5827

//MAC_4528 replaced by MAC_5827

//MAC_4527 replaced by MAC_5826

//MAC_4526 replaced by MAC_5827

//MAC_4525 replaced by MAC_5827

//MAC_4524 replaced by MAC_5826

//MAC_4535 replaced by MAC_5827

//MAC_4534 replaced by MAC_5827

//MAC_4533 replaced by MAC_5826

//MAC_4532 replaced by MAC_5827

//MAC_4531 replaced by MAC_5827

//MAC_4530 replaced by MAC_5826

//MAC_4541 replaced by MAC_5827

//MAC_4540 replaced by MAC_5827

//MAC_4539 replaced by MAC_5826

//MAC_4538 replaced by MAC_5827

//MAC_4537 replaced by MAC_5827

//MAC_4536 replaced by MAC_5826

//MAC_4547 replaced by MAC_5827

//MAC_4546 replaced by MAC_5827

//MAC_4545 replaced by MAC_5826

//MAC_4544 replaced by MAC_5827

//MAC_4543 replaced by MAC_5827

//MAC_4542 replaced by MAC_5826

//MAC_4553 replaced by MAC_5827

//MAC_4552 replaced by MAC_5827

//MAC_4551 replaced by MAC_5826

//MAC_4550 replaced by MAC_5827

//MAC_4549 replaced by MAC_5827

//MAC_4548 replaced by MAC_5826

//MAC_4559 replaced by MAC_5827

//MAC_4558 replaced by MAC_5827

//MAC_4557 replaced by MAC_5826

//MAC_4556 replaced by MAC_5827

//MAC_4555 replaced by MAC_5827

//MAC_4554 replaced by MAC_5826

//MAC_4565 replaced by MAC_5827

//MAC_4564 replaced by MAC_5827

//MAC_4563 replaced by MAC_5826

//MAC_4562 replaced by MAC_5827

//MAC_4561 replaced by MAC_5827

//MAC_4560 replaced by MAC_5826

//MAC_4571 replaced by MAC_5827

//MAC_4570 replaced by MAC_5827

//MAC_4569 replaced by MAC_5826

//MAC_4568 replaced by MAC_5827

//MAC_4567 replaced by MAC_5827

//MAC_4566 replaced by MAC_5826

//MAC_4577 replaced by MAC_5827

//MAC_4576 replaced by MAC_5827

//MAC_4575 replaced by MAC_5826

//MAC_4574 replaced by MAC_5827

//MAC_4573 replaced by MAC_5827

//MAC_4572 replaced by MAC_5826

//MAC_4583 replaced by MAC_5827

//MAC_4582 replaced by MAC_5827

//MAC_4581 replaced by MAC_5826

//MAC_4580 replaced by MAC_5827

//MAC_4579 replaced by MAC_5827

//MAC_4578 replaced by MAC_5826

//MAC_4589 replaced by MAC_5827

//MAC_4588 replaced by MAC_5827

//MAC_4587 replaced by MAC_5826

//MAC_4586 replaced by MAC_5827

//MAC_4585 replaced by MAC_5827

//MAC_4584 replaced by MAC_5826

//MAC_4595 replaced by MAC_5827

//MAC_4594 replaced by MAC_5827

//MAC_4593 replaced by MAC_5826

//MAC_4592 replaced by MAC_5827

//MAC_4591 replaced by MAC_5827

//MAC_4590 replaced by MAC_5826

//MAC_4601 replaced by MAC_5827

//MAC_4600 replaced by MAC_5827

//MAC_4599 replaced by MAC_5826

//MAC_4598 replaced by MAC_5827

//MAC_4597 replaced by MAC_5827

//MAC_4596 replaced by MAC_5826

//MAC_4607 replaced by MAC_5827

//MAC_4606 replaced by MAC_5827

//MAC_4605 replaced by MAC_5826

//MAC_4604 replaced by MAC_5827

//MAC_4603 replaced by MAC_5827

//MAC_4602 replaced by MAC_5826

//MAC_4613 replaced by MAC_5827

//MAC_4612 replaced by MAC_5827

//MAC_4611 replaced by MAC_5826

//MAC_4610 replaced by MAC_5827

//MAC_4609 replaced by MAC_5827

//MAC_4608 replaced by MAC_5826

//MAC_4619 replaced by MAC_5827

//MAC_4618 replaced by MAC_5827

//MAC_4617 replaced by MAC_5826

//MAC_4616 replaced by MAC_5827

//MAC_4615 replaced by MAC_5827

//MAC_4614 replaced by MAC_5826

//MAC_4625 replaced by MAC_5827

//MAC_4624 replaced by MAC_5827

//MAC_4623 replaced by MAC_5826

//MAC_4622 replaced by MAC_5827

//MAC_4621 replaced by MAC_5827

//MAC_4620 replaced by MAC_5826

//MAC_4631 replaced by MAC_5827

//MAC_4630 replaced by MAC_5827

//MAC_4629 replaced by MAC_5826

//MAC_4628 replaced by MAC_5827

//MAC_4627 replaced by MAC_5827

//MAC_4626 replaced by MAC_5826

//MAC_4637 replaced by MAC_5827

//MAC_4636 replaced by MAC_5827

//MAC_4635 replaced by MAC_5826

//MAC_4634 replaced by MAC_5827

//MAC_4633 replaced by MAC_5827

//MAC_4632 replaced by MAC_5826

//MAC_4643 replaced by MAC_5827

//MAC_4642 replaced by MAC_5827

//MAC_4641 replaced by MAC_5826

//MAC_4640 replaced by MAC_5827

//MAC_4639 replaced by MAC_5827

//MAC_4638 replaced by MAC_5826

//MAC_4649 replaced by MAC_5827

//MAC_4648 replaced by MAC_5827

//MAC_4647 replaced by MAC_5826

//MAC_4646 replaced by MAC_5827

//MAC_4645 replaced by MAC_5827

//MAC_4644 replaced by MAC_5826

//MAC_4655 replaced by MAC_5827

//MAC_4654 replaced by MAC_5827

//MAC_4653 replaced by MAC_5826

//MAC_4652 replaced by MAC_5827

//MAC_4651 replaced by MAC_5827

//MAC_4650 replaced by MAC_5826

//MAC_4661 replaced by MAC_5827

//MAC_4660 replaced by MAC_5827

//MAC_4659 replaced by MAC_5826

//MAC_4658 replaced by MAC_5827

//MAC_4657 replaced by MAC_5827

//MAC_4656 replaced by MAC_5826

//MAC_4667 replaced by MAC_5827

//MAC_4666 replaced by MAC_5827

//MAC_4665 replaced by MAC_5826

//MAC_4664 replaced by MAC_5827

//MAC_4663 replaced by MAC_5827

//MAC_4662 replaced by MAC_5826

//MAC_4673 replaced by MAC_5827

//MAC_4672 replaced by MAC_5827

//MAC_4671 replaced by MAC_5826

//MAC_4670 replaced by MAC_5827

//MAC_4669 replaced by MAC_5827

//MAC_4668 replaced by MAC_5826

//MAC_4679 replaced by MAC_5827

//MAC_4678 replaced by MAC_5827

//MAC_4677 replaced by MAC_5826

//MAC_4676 replaced by MAC_5827

//MAC_4675 replaced by MAC_5827

//MAC_4674 replaced by MAC_5826

//MAC_4685 replaced by MAC_5827

//MAC_4684 replaced by MAC_5827

//MAC_4683 replaced by MAC_5826

//MAC_4682 replaced by MAC_5827

//MAC_4681 replaced by MAC_5827

//MAC_4680 replaced by MAC_5826

//MAC_4691 replaced by MAC_5827

//MAC_4690 replaced by MAC_5827

//MAC_4689 replaced by MAC_5826

//MAC_4688 replaced by MAC_5827

//MAC_4687 replaced by MAC_5827

//MAC_4686 replaced by MAC_5826

//MAC_4697 replaced by MAC_5827

//MAC_4696 replaced by MAC_5827

//MAC_4695 replaced by MAC_5826

//MAC_4694 replaced by MAC_5827

//MAC_4693 replaced by MAC_5827

//MAC_4692 replaced by MAC_5826

//MAC_4703 replaced by MAC_5827

//MAC_4702 replaced by MAC_5827

//MAC_4701 replaced by MAC_5826

//MAC_4700 replaced by MAC_5827

//MAC_4699 replaced by MAC_5827

//MAC_4698 replaced by MAC_5826

//MAC_4709 replaced by MAC_5827

//MAC_4708 replaced by MAC_5827

//MAC_4707 replaced by MAC_5826

//MAC_4706 replaced by MAC_5827

//MAC_4705 replaced by MAC_5827

//MAC_4704 replaced by MAC_5826

//MAC_4715 replaced by MAC_5827

//MAC_4714 replaced by MAC_5827

//MAC_4713 replaced by MAC_5826

//MAC_4712 replaced by MAC_5827

//MAC_4711 replaced by MAC_5827

//MAC_4710 replaced by MAC_5826

//MAC_4721 replaced by MAC_5827

//MAC_4720 replaced by MAC_5827

//MAC_4719 replaced by MAC_5826

//MAC_4718 replaced by MAC_5827

//MAC_4717 replaced by MAC_5827

//MAC_4716 replaced by MAC_5826

//MAC_4727 replaced by MAC_5827

//MAC_4726 replaced by MAC_5827

//MAC_4725 replaced by MAC_5826

//MAC_4724 replaced by MAC_5827

//MAC_4723 replaced by MAC_5827

//MAC_4722 replaced by MAC_5826

//MAC_4733 replaced by MAC_5827

//MAC_4732 replaced by MAC_5827

//MAC_4731 replaced by MAC_5826

//MAC_4730 replaced by MAC_5827

//MAC_4729 replaced by MAC_5827

//MAC_4728 replaced by MAC_5826

//MAC_4739 replaced by MAC_5827

//MAC_4738 replaced by MAC_5827

//MAC_4737 replaced by MAC_5826

//MAC_4736 replaced by MAC_5827

//MAC_4735 replaced by MAC_5827

//MAC_4734 replaced by MAC_5826

//MAC_4745 replaced by MAC_5827

//MAC_4744 replaced by MAC_5827

//MAC_4743 replaced by MAC_5826

//MAC_4742 replaced by MAC_5827

//MAC_4741 replaced by MAC_5827

//MAC_4740 replaced by MAC_5826

//MAC_4751 replaced by MAC_5827

//MAC_4750 replaced by MAC_5827

//MAC_4749 replaced by MAC_5826

//MAC_4748 replaced by MAC_5827

//MAC_4747 replaced by MAC_5827

//MAC_4746 replaced by MAC_5826

//MAC_4757 replaced by MAC_5827

//MAC_4756 replaced by MAC_5827

//MAC_4755 replaced by MAC_5826

//MAC_4754 replaced by MAC_5827

//MAC_4753 replaced by MAC_5827

//MAC_4752 replaced by MAC_5826

//MAC_4763 replaced by MAC_5827

//MAC_4762 replaced by MAC_5827

//MAC_4761 replaced by MAC_5826

//MAC_4760 replaced by MAC_5827

//MAC_4759 replaced by MAC_5827

//MAC_4758 replaced by MAC_5826

//MAC_4769 replaced by MAC_5827

//MAC_4768 replaced by MAC_5827

//MAC_4767 replaced by MAC_5826

//MAC_4766 replaced by MAC_5827

//MAC_4765 replaced by MAC_5827

//MAC_4764 replaced by MAC_5826

//MAC_4775 replaced by MAC_5827

//MAC_4774 replaced by MAC_5827

//MAC_4773 replaced by MAC_5826

//MAC_4772 replaced by MAC_5827

//MAC_4771 replaced by MAC_5827

//MAC_4770 replaced by MAC_5826

//MAC_4781 replaced by MAC_5827

//MAC_4780 replaced by MAC_5827

//MAC_4779 replaced by MAC_5826

//MAC_4778 replaced by MAC_5827

//MAC_4777 replaced by MAC_5827

//MAC_4776 replaced by MAC_5826

//MAC_4787 replaced by MAC_5827

//MAC_4786 replaced by MAC_5827

//MAC_4785 replaced by MAC_5826

//MAC_4784 replaced by MAC_5827

//MAC_4783 replaced by MAC_5827

//MAC_4782 replaced by MAC_5826

//MAC_4793 replaced by MAC_5827

//MAC_4792 replaced by MAC_5827

//MAC_4791 replaced by MAC_5826

//MAC_4790 replaced by MAC_5827

//MAC_4789 replaced by MAC_5827

//MAC_4788 replaced by MAC_5826

//MAC_4799 replaced by MAC_5827

//MAC_4798 replaced by MAC_5827

//MAC_4797 replaced by MAC_5826

//MAC_4796 replaced by MAC_5827

//MAC_4795 replaced by MAC_5827

//MAC_4794 replaced by MAC_5826

//MAC_4805 replaced by MAC_5827

//MAC_4804 replaced by MAC_5827

//MAC_4803 replaced by MAC_5826

//MAC_4802 replaced by MAC_5827

//MAC_4801 replaced by MAC_5827

//MAC_4800 replaced by MAC_5826

//MAC_4811 replaced by MAC_5827

//MAC_4810 replaced by MAC_5827

//MAC_4809 replaced by MAC_5826

//MAC_4808 replaced by MAC_5827

//MAC_4807 replaced by MAC_5827

//MAC_4806 replaced by MAC_5826

//MAC_4817 replaced by MAC_5827

//MAC_4816 replaced by MAC_5827

//MAC_4815 replaced by MAC_5826

//MAC_4814 replaced by MAC_5827

//MAC_4813 replaced by MAC_5827

//MAC_4812 replaced by MAC_5826

//MAC_4823 replaced by MAC_5827

//MAC_4822 replaced by MAC_5827

//MAC_4821 replaced by MAC_5826

//MAC_4820 replaced by MAC_5827

//MAC_4819 replaced by MAC_5827

//MAC_4818 replaced by MAC_5826

//MAC_4829 replaced by MAC_5827

//MAC_4828 replaced by MAC_5827

//MAC_4827 replaced by MAC_5826

//MAC_4826 replaced by MAC_5827

//MAC_4825 replaced by MAC_5827

//MAC_4824 replaced by MAC_5826

//MAC_4835 replaced by MAC_5827

//MAC_4834 replaced by MAC_5827

//MAC_4833 replaced by MAC_5826

//MAC_4832 replaced by MAC_5827

//MAC_4831 replaced by MAC_5827

//MAC_4830 replaced by MAC_5826

//MAC_4841 replaced by MAC_5827

//MAC_4840 replaced by MAC_5827

//MAC_4839 replaced by MAC_5826

//MAC_4838 replaced by MAC_5827

//MAC_4837 replaced by MAC_5827

//MAC_4836 replaced by MAC_5826

//MAC_4847 replaced by MAC_5827

//MAC_4846 replaced by MAC_5827

//MAC_4845 replaced by MAC_5826

//MAC_4844 replaced by MAC_5827

//MAC_4843 replaced by MAC_5827

//MAC_4842 replaced by MAC_5826

//MAC_4853 replaced by MAC_5827

//MAC_4852 replaced by MAC_5827

//MAC_4851 replaced by MAC_5826

//MAC_4850 replaced by MAC_5827

//MAC_4849 replaced by MAC_5827

//MAC_4848 replaced by MAC_5826

//MAC_4859 replaced by MAC_5827

//MAC_4858 replaced by MAC_5827

//MAC_4857 replaced by MAC_5826

//MAC_4856 replaced by MAC_5827

//MAC_4855 replaced by MAC_5827

//MAC_4854 replaced by MAC_5826

//MAC_4865 replaced by MAC_5827

//MAC_4864 replaced by MAC_5827

//MAC_4863 replaced by MAC_5826

//MAC_4862 replaced by MAC_5827

//MAC_4861 replaced by MAC_5827

//MAC_4860 replaced by MAC_5826

//MAC_4871 replaced by MAC_5827

//MAC_4870 replaced by MAC_5827

//MAC_4869 replaced by MAC_5826

//MAC_4868 replaced by MAC_5827

//MAC_4867 replaced by MAC_5827

//MAC_4866 replaced by MAC_5826

//MAC_4877 replaced by MAC_5827

//MAC_4876 replaced by MAC_5827

//MAC_4875 replaced by MAC_5826

//MAC_4874 replaced by MAC_5827

//MAC_4873 replaced by MAC_5827

//MAC_4872 replaced by MAC_5826

//MAC_4883 replaced by MAC_5827

//MAC_4882 replaced by MAC_5827

//MAC_4881 replaced by MAC_5826

//MAC_4880 replaced by MAC_5827

//MAC_4879 replaced by MAC_5827

//MAC_4878 replaced by MAC_5826

//MAC_4889 replaced by MAC_5827

//MAC_4888 replaced by MAC_5827

//MAC_4887 replaced by MAC_5826

//MAC_4886 replaced by MAC_5827

//MAC_4885 replaced by MAC_5827

//MAC_4884 replaced by MAC_5826

//MAC_4895 replaced by MAC_5827

//MAC_4894 replaced by MAC_5827

//MAC_4893 replaced by MAC_5826

//MAC_4892 replaced by MAC_5827

//MAC_4891 replaced by MAC_5827

//MAC_4890 replaced by MAC_5826

//MAC_4901 replaced by MAC_5827

//MAC_4900 replaced by MAC_5827

//MAC_4899 replaced by MAC_5826

//MAC_4898 replaced by MAC_5827

//MAC_4897 replaced by MAC_5827

//MAC_4896 replaced by MAC_5826

//MAC_4907 replaced by MAC_5827

//MAC_4906 replaced by MAC_5827

//MAC_4905 replaced by MAC_5826

//MAC_4904 replaced by MAC_5827

//MAC_4903 replaced by MAC_5827

//MAC_4902 replaced by MAC_5826

//MAC_4913 replaced by MAC_5827

//MAC_4912 replaced by MAC_5827

//MAC_4911 replaced by MAC_5826

//MAC_4910 replaced by MAC_5827

//MAC_4909 replaced by MAC_5827

//MAC_4908 replaced by MAC_5826

//MAC_4919 replaced by MAC_5827

//MAC_4918 replaced by MAC_5827

//MAC_4917 replaced by MAC_5826

//MAC_4916 replaced by MAC_5827

//MAC_4915 replaced by MAC_5827

//MAC_4914 replaced by MAC_5826

//MAC_4925 replaced by MAC_5827

//MAC_4924 replaced by MAC_5827

//MAC_4923 replaced by MAC_5826

//MAC_4922 replaced by MAC_5827

//MAC_4921 replaced by MAC_5827

//MAC_4920 replaced by MAC_5826

//MAC_4931 replaced by MAC_5827

//MAC_4930 replaced by MAC_5827

//MAC_4929 replaced by MAC_5826

//MAC_4928 replaced by MAC_5827

//MAC_4927 replaced by MAC_5827

//MAC_4926 replaced by MAC_5826

//MAC_4937 replaced by MAC_5827

//MAC_4936 replaced by MAC_5827

//MAC_4935 replaced by MAC_5826

//MAC_4934 replaced by MAC_5827

//MAC_4933 replaced by MAC_5827

//MAC_4932 replaced by MAC_5826

//MAC_4943 replaced by MAC_5827

//MAC_4942 replaced by MAC_5827

//MAC_4941 replaced by MAC_5826

//MAC_4940 replaced by MAC_5827

//MAC_4939 replaced by MAC_5827

//MAC_4938 replaced by MAC_5826

//MAC_4949 replaced by MAC_5827

//MAC_4948 replaced by MAC_5827

//MAC_4947 replaced by MAC_5826

//MAC_4946 replaced by MAC_5827

//MAC_4945 replaced by MAC_5827

//MAC_4944 replaced by MAC_5826

//MAC_4955 replaced by MAC_5827

//MAC_4954 replaced by MAC_5827

//MAC_4953 replaced by MAC_5826

//MAC_4952 replaced by MAC_5827

//MAC_4951 replaced by MAC_5827

//MAC_4950 replaced by MAC_5826

//MAC_4961 replaced by MAC_5827

//MAC_4960 replaced by MAC_5827

//MAC_4959 replaced by MAC_5826

//MAC_4958 replaced by MAC_5827

//MAC_4957 replaced by MAC_5827

//MAC_4956 replaced by MAC_5826

//MAC_4967 replaced by MAC_5827

//MAC_4966 replaced by MAC_5827

//MAC_4965 replaced by MAC_5826

//MAC_4964 replaced by MAC_5827

//MAC_4963 replaced by MAC_5827

//MAC_4962 replaced by MAC_5826

//MAC_4973 replaced by MAC_5827

//MAC_4972 replaced by MAC_5827

//MAC_4971 replaced by MAC_5826

//MAC_4970 replaced by MAC_5827

//MAC_4969 replaced by MAC_5827

//MAC_4968 replaced by MAC_5826

//MAC_4979 replaced by MAC_5827

//MAC_4978 replaced by MAC_5827

//MAC_4977 replaced by MAC_5826

//MAC_4976 replaced by MAC_5827

//MAC_4975 replaced by MAC_5827

//MAC_4974 replaced by MAC_5826

//MAC_4985 replaced by MAC_5827

//MAC_4984 replaced by MAC_5827

//MAC_4983 replaced by MAC_5826

//MAC_4982 replaced by MAC_5827

//MAC_4981 replaced by MAC_5827

//MAC_4980 replaced by MAC_5826

//MAC_4991 replaced by MAC_5827

//MAC_4990 replaced by MAC_5827

//MAC_4989 replaced by MAC_5826

//MAC_4988 replaced by MAC_5827

//MAC_4987 replaced by MAC_5827

//MAC_4986 replaced by MAC_5826

//MAC_4997 replaced by MAC_5827

//MAC_4996 replaced by MAC_5827

//MAC_4995 replaced by MAC_5826

//MAC_4994 replaced by MAC_5827

//MAC_4993 replaced by MAC_5827

//MAC_4992 replaced by MAC_5826

//MAC_5003 replaced by MAC_5827

//MAC_5002 replaced by MAC_5827

//MAC_5001 replaced by MAC_5826

//MAC_5000 replaced by MAC_5827

//MAC_4999 replaced by MAC_5827

//MAC_4998 replaced by MAC_5826

//MAC_5009 replaced by MAC_5827

//MAC_5008 replaced by MAC_5827

//MAC_5007 replaced by MAC_5826

//MAC_5006 replaced by MAC_5827

//MAC_5005 replaced by MAC_5827

//MAC_5004 replaced by MAC_5826

//MAC_5015 replaced by MAC_5827

//MAC_5014 replaced by MAC_5827

//MAC_5013 replaced by MAC_5826

//MAC_5012 replaced by MAC_5827

//MAC_5011 replaced by MAC_5827

//MAC_5010 replaced by MAC_5826

//MAC_5021 replaced by MAC_5827

//MAC_5020 replaced by MAC_5827

//MAC_5019 replaced by MAC_5826

//MAC_5018 replaced by MAC_5827

//MAC_5017 replaced by MAC_5827

//MAC_5016 replaced by MAC_5826

//MAC_5027 replaced by MAC_5827

//MAC_5026 replaced by MAC_5827

//MAC_5025 replaced by MAC_5826

//MAC_5024 replaced by MAC_5827

//MAC_5023 replaced by MAC_5827

//MAC_5022 replaced by MAC_5826

//MAC_5033 replaced by MAC_5827

//MAC_5032 replaced by MAC_5827

//MAC_5031 replaced by MAC_5826

//MAC_5030 replaced by MAC_5827

//MAC_5029 replaced by MAC_5827

//MAC_5028 replaced by MAC_5826

//MAC_5039 replaced by MAC_5827

//MAC_5038 replaced by MAC_5827

//MAC_5037 replaced by MAC_5826

//MAC_5036 replaced by MAC_5827

//MAC_5035 replaced by MAC_5827

//MAC_5034 replaced by MAC_5826

//MAC_5045 replaced by MAC_5827

//MAC_5044 replaced by MAC_5827

//MAC_5043 replaced by MAC_5826

//MAC_5042 replaced by MAC_5827

//MAC_5041 replaced by MAC_5827

//MAC_5040 replaced by MAC_5826

//MAC_5051 replaced by MAC_5827

//MAC_5050 replaced by MAC_5827

//MAC_5049 replaced by MAC_5826

//MAC_5048 replaced by MAC_5827

//MAC_5047 replaced by MAC_5827

//MAC_5046 replaced by MAC_5826

//MAC_5057 replaced by MAC_5827

//MAC_5056 replaced by MAC_5827

//MAC_5055 replaced by MAC_5826

//MAC_5054 replaced by MAC_5827

//MAC_5053 replaced by MAC_5827

//MAC_5052 replaced by MAC_5826

//MAC_5063 replaced by MAC_5827

//MAC_5062 replaced by MAC_5827

//MAC_5061 replaced by MAC_5826

//MAC_5060 replaced by MAC_5827

//MAC_5059 replaced by MAC_5827

//MAC_5058 replaced by MAC_5826

//MAC_5069 replaced by MAC_5827

//MAC_5068 replaced by MAC_5827

//MAC_5067 replaced by MAC_5826

//MAC_5066 replaced by MAC_5827

//MAC_5065 replaced by MAC_5827

//MAC_5064 replaced by MAC_5826

//MAC_5075 replaced by MAC_5827

//MAC_5074 replaced by MAC_5827

//MAC_5073 replaced by MAC_5826

//MAC_5072 replaced by MAC_5827

//MAC_5071 replaced by MAC_5827

//MAC_5070 replaced by MAC_5826

//MAC_5081 replaced by MAC_5827

//MAC_5080 replaced by MAC_5827

//MAC_5079 replaced by MAC_5826

//MAC_5078 replaced by MAC_5827

//MAC_5077 replaced by MAC_5827

//MAC_5076 replaced by MAC_5826

//MAC_5087 replaced by MAC_5827

//MAC_5086 replaced by MAC_5827

//MAC_5085 replaced by MAC_5826

//MAC_5084 replaced by MAC_5827

//MAC_5083 replaced by MAC_5827

//MAC_5082 replaced by MAC_5826

//MAC_5093 replaced by MAC_5827

//MAC_5092 replaced by MAC_5827

//MAC_5091 replaced by MAC_5826

//MAC_5090 replaced by MAC_5827

//MAC_5089 replaced by MAC_5827

//MAC_5088 replaced by MAC_5826

//MAC_5099 replaced by MAC_5827

//MAC_5098 replaced by MAC_5827

//MAC_5097 replaced by MAC_5826

//MAC_5096 replaced by MAC_5827

//MAC_5095 replaced by MAC_5827

//MAC_5094 replaced by MAC_5826

//MAC_5105 replaced by MAC_5827

//MAC_5104 replaced by MAC_5827

//MAC_5103 replaced by MAC_5826

//MAC_5102 replaced by MAC_5827

//MAC_5101 replaced by MAC_5827

//MAC_5100 replaced by MAC_5826

//MAC_5111 replaced by MAC_5827

//MAC_5110 replaced by MAC_5827

//MAC_5109 replaced by MAC_5826

//MAC_5108 replaced by MAC_5827

//MAC_5107 replaced by MAC_5827

//MAC_5106 replaced by MAC_5826

//MAC_5117 replaced by MAC_5827

//MAC_5116 replaced by MAC_5827

//MAC_5115 replaced by MAC_5826

//MAC_5114 replaced by MAC_5827

//MAC_5113 replaced by MAC_5827

//MAC_5112 replaced by MAC_5826

//MAC_5123 replaced by MAC_5827

//MAC_5122 replaced by MAC_5827

//MAC_5121 replaced by MAC_5826

//MAC_5120 replaced by MAC_5827

//MAC_5119 replaced by MAC_5827

//MAC_5118 replaced by MAC_5826

//MAC_5129 replaced by MAC_5827

//MAC_5128 replaced by MAC_5827

//MAC_5127 replaced by MAC_5826

//MAC_5126 replaced by MAC_5827

//MAC_5125 replaced by MAC_5827

//MAC_5124 replaced by MAC_5826

//MAC_5135 replaced by MAC_5827

//MAC_5134 replaced by MAC_5827

//MAC_5133 replaced by MAC_5826

//MAC_5132 replaced by MAC_5827

//MAC_5131 replaced by MAC_5827

//MAC_5130 replaced by MAC_5826

//MAC_5141 replaced by MAC_5827

//MAC_5140 replaced by MAC_5827

//MAC_5139 replaced by MAC_5826

//MAC_5138 replaced by MAC_5827

//MAC_5137 replaced by MAC_5827

//MAC_5136 replaced by MAC_5826

//MAC_5147 replaced by MAC_5827

//MAC_5146 replaced by MAC_5827

//MAC_5145 replaced by MAC_5826

//MAC_5144 replaced by MAC_5827

//MAC_5143 replaced by MAC_5827

//MAC_5142 replaced by MAC_5826

//MAC_5153 replaced by MAC_5827

//MAC_5152 replaced by MAC_5827

//MAC_5151 replaced by MAC_5826

//MAC_5150 replaced by MAC_5827

//MAC_5149 replaced by MAC_5827

//MAC_5148 replaced by MAC_5826

//MAC_5159 replaced by MAC_5827

//MAC_5158 replaced by MAC_5827

//MAC_5157 replaced by MAC_5826

//MAC_5156 replaced by MAC_5827

//MAC_5155 replaced by MAC_5827

//MAC_5154 replaced by MAC_5826

//MAC_5165 replaced by MAC_5827

//MAC_5164 replaced by MAC_5827

//MAC_5163 replaced by MAC_5826

//MAC_5162 replaced by MAC_5827

//MAC_5161 replaced by MAC_5827

//MAC_5160 replaced by MAC_5826

//MAC_5171 replaced by MAC_5827

//MAC_5170 replaced by MAC_5827

//MAC_5169 replaced by MAC_5826

//MAC_5168 replaced by MAC_5827

//MAC_5167 replaced by MAC_5827

//MAC_5166 replaced by MAC_5826

//MAC_5177 replaced by MAC_5827

//MAC_5176 replaced by MAC_5827

//MAC_5175 replaced by MAC_5826

//MAC_5174 replaced by MAC_5827

//MAC_5173 replaced by MAC_5827

//MAC_5172 replaced by MAC_5826

//MAC_5183 replaced by MAC_5827

//MAC_5182 replaced by MAC_5827

//MAC_5181 replaced by MAC_5826

//MAC_5180 replaced by MAC_5827

//MAC_5179 replaced by MAC_5827

//MAC_5178 replaced by MAC_5826

//MAC_5189 replaced by MAC_5827

//MAC_5188 replaced by MAC_5827

//MAC_5187 replaced by MAC_5826

//MAC_5186 replaced by MAC_5827

//MAC_5185 replaced by MAC_5827

//MAC_5184 replaced by MAC_5826

//MAC_5195 replaced by MAC_5827

//MAC_5194 replaced by MAC_5827

//MAC_5193 replaced by MAC_5826

//MAC_5192 replaced by MAC_5827

//MAC_5191 replaced by MAC_5827

//MAC_5190 replaced by MAC_5826

//MAC_5201 replaced by MAC_5827

//MAC_5200 replaced by MAC_5827

//MAC_5199 replaced by MAC_5826

//MAC_5198 replaced by MAC_5827

//MAC_5197 replaced by MAC_5827

//MAC_5196 replaced by MAC_5826

//MAC_5207 replaced by MAC_5827

//MAC_5206 replaced by MAC_5827

//MAC_5205 replaced by MAC_5826

//MAC_5204 replaced by MAC_5827

//MAC_5203 replaced by MAC_5827

//MAC_5202 replaced by MAC_5826

//MAC_5213 replaced by MAC_5827

//MAC_5212 replaced by MAC_5827

//MAC_5211 replaced by MAC_5826

//MAC_5210 replaced by MAC_5827

//MAC_5209 replaced by MAC_5827

//MAC_5208 replaced by MAC_5826

//MAC_5219 replaced by MAC_5827

//MAC_5218 replaced by MAC_5827

//MAC_5217 replaced by MAC_5826

//MAC_5216 replaced by MAC_5827

//MAC_5215 replaced by MAC_5827

//MAC_5214 replaced by MAC_5826

//MAC_5225 replaced by MAC_5827

//MAC_5224 replaced by MAC_5827

//MAC_5223 replaced by MAC_5826

//MAC_5222 replaced by MAC_5827

//MAC_5221 replaced by MAC_5827

//MAC_5220 replaced by MAC_5826

//MAC_5231 replaced by MAC_5827

//MAC_5230 replaced by MAC_5827

//MAC_5229 replaced by MAC_5826

//MAC_5228 replaced by MAC_5827

//MAC_5227 replaced by MAC_5827

//MAC_5226 replaced by MAC_5826

//MAC_5237 replaced by MAC_5827

//MAC_5236 replaced by MAC_5827

//MAC_5235 replaced by MAC_5826

//MAC_5234 replaced by MAC_5827

//MAC_5233 replaced by MAC_5827

//MAC_5232 replaced by MAC_5826

//MAC_5243 replaced by MAC_5827

//MAC_5242 replaced by MAC_5827

//MAC_5241 replaced by MAC_5826

//MAC_5240 replaced by MAC_5827

//MAC_5239 replaced by MAC_5827

//MAC_5238 replaced by MAC_5826

//MAC_5249 replaced by MAC_5827

//MAC_5248 replaced by MAC_5827

//MAC_5247 replaced by MAC_5826

//MAC_5246 replaced by MAC_5827

//MAC_5245 replaced by MAC_5827

//MAC_5244 replaced by MAC_5826

//MAC_5255 replaced by MAC_5827

//MAC_5254 replaced by MAC_5827

//MAC_5253 replaced by MAC_5826

//MAC_5252 replaced by MAC_5827

//MAC_5251 replaced by MAC_5827

//MAC_5250 replaced by MAC_5826

//MAC_5261 replaced by MAC_5827

//MAC_5260 replaced by MAC_5827

//MAC_5259 replaced by MAC_5826

//MAC_5258 replaced by MAC_5827

//MAC_5257 replaced by MAC_5827

//MAC_5256 replaced by MAC_5826

//MAC_5267 replaced by MAC_5827

//MAC_5266 replaced by MAC_5827

//MAC_5265 replaced by MAC_5826

//MAC_5264 replaced by MAC_5827

//MAC_5263 replaced by MAC_5827

//MAC_5262 replaced by MAC_5826

//MAC_5273 replaced by MAC_5827

//MAC_5272 replaced by MAC_5827

//MAC_5271 replaced by MAC_5826

//MAC_5270 replaced by MAC_5827

//MAC_5269 replaced by MAC_5827

//MAC_5268 replaced by MAC_5826

//MAC_5279 replaced by MAC_5827

//MAC_5278 replaced by MAC_5827

//MAC_5277 replaced by MAC_5826

//MAC_5276 replaced by MAC_5827

//MAC_5275 replaced by MAC_5827

//MAC_5274 replaced by MAC_5826

//MAC_5285 replaced by MAC_5827

//MAC_5284 replaced by MAC_5827

//MAC_5283 replaced by MAC_5826

//MAC_5282 replaced by MAC_5827

//MAC_5281 replaced by MAC_5827

//MAC_5280 replaced by MAC_5826

//MAC_5291 replaced by MAC_5827

//MAC_5290 replaced by MAC_5827

//MAC_5289 replaced by MAC_5826

//MAC_5288 replaced by MAC_5827

//MAC_5287 replaced by MAC_5827

//MAC_5286 replaced by MAC_5826

//MAC_5297 replaced by MAC_5827

//MAC_5296 replaced by MAC_5827

//MAC_5295 replaced by MAC_5826

//MAC_5294 replaced by MAC_5827

//MAC_5293 replaced by MAC_5827

//MAC_5292 replaced by MAC_5826

//MAC_5303 replaced by MAC_5827

//MAC_5302 replaced by MAC_5827

//MAC_5301 replaced by MAC_5826

//MAC_5300 replaced by MAC_5827

//MAC_5299 replaced by MAC_5827

//MAC_5298 replaced by MAC_5826

//MAC_5309 replaced by MAC_5827

//MAC_5308 replaced by MAC_5827

//MAC_5307 replaced by MAC_5826

//MAC_5306 replaced by MAC_5827

//MAC_5305 replaced by MAC_5827

//MAC_5304 replaced by MAC_5826

//MAC_5315 replaced by MAC_5827

//MAC_5314 replaced by MAC_5827

//MAC_5313 replaced by MAC_5826

//MAC_5312 replaced by MAC_5827

//MAC_5311 replaced by MAC_5827

//MAC_5310 replaced by MAC_5826

//MAC_5321 replaced by MAC_5827

//MAC_5320 replaced by MAC_5827

//MAC_5319 replaced by MAC_5826

//MAC_5318 replaced by MAC_5827

//MAC_5317 replaced by MAC_5827

//MAC_5316 replaced by MAC_5826

//MAC_5327 replaced by MAC_5827

//MAC_5326 replaced by MAC_5827

//MAC_5325 replaced by MAC_5826

//MAC_5324 replaced by MAC_5827

//MAC_5323 replaced by MAC_5827

//MAC_5322 replaced by MAC_5826

//MAC_5333 replaced by MAC_5827

//MAC_5332 replaced by MAC_5827

//MAC_5331 replaced by MAC_5826

//MAC_5330 replaced by MAC_5827

//MAC_5329 replaced by MAC_5827

//MAC_5328 replaced by MAC_5826

//MAC_5339 replaced by MAC_5827

//MAC_5338 replaced by MAC_5827

//MAC_5337 replaced by MAC_5826

//MAC_5336 replaced by MAC_5827

//MAC_5335 replaced by MAC_5827

//MAC_5334 replaced by MAC_5826

//MAC_5345 replaced by MAC_5827

//MAC_5344 replaced by MAC_5827

//MAC_5343 replaced by MAC_5826

//MAC_5342 replaced by MAC_5827

//MAC_5341 replaced by MAC_5827

//MAC_5340 replaced by MAC_5826

//MAC_5351 replaced by MAC_5827

//MAC_5350 replaced by MAC_5827

//MAC_5349 replaced by MAC_5826

//MAC_5348 replaced by MAC_5827

//MAC_5347 replaced by MAC_5827

//MAC_5346 replaced by MAC_5826

//MAC_5357 replaced by MAC_5827

//MAC_5356 replaced by MAC_5827

//MAC_5355 replaced by MAC_5826

//MAC_5354 replaced by MAC_5827

//MAC_5353 replaced by MAC_5827

//MAC_5352 replaced by MAC_5826

//MAC_5363 replaced by MAC_5827

//MAC_5362 replaced by MAC_5827

//MAC_5361 replaced by MAC_5826

//MAC_5360 replaced by MAC_5827

//MAC_5359 replaced by MAC_5827

//MAC_5358 replaced by MAC_5826

//MAC_5369 replaced by MAC_5827

//MAC_5368 replaced by MAC_5827

//MAC_5367 replaced by MAC_5826

//MAC_5366 replaced by MAC_5827

//MAC_5365 replaced by MAC_5827

//MAC_5364 replaced by MAC_5826

//MAC_5375 replaced by MAC_5827

//MAC_5374 replaced by MAC_5827

//MAC_5373 replaced by MAC_5826

//MAC_5372 replaced by MAC_5827

//MAC_5371 replaced by MAC_5827

//MAC_5370 replaced by MAC_5826

//MAC_5381 replaced by MAC_5827

//MAC_5380 replaced by MAC_5827

//MAC_5379 replaced by MAC_5826

//MAC_5378 replaced by MAC_5827

//MAC_5377 replaced by MAC_5827

//MAC_5376 replaced by MAC_5826

//MAC_5387 replaced by MAC_5827

//MAC_5386 replaced by MAC_5827

//MAC_5385 replaced by MAC_5826

//MAC_5384 replaced by MAC_5827

//MAC_5383 replaced by MAC_5827

//MAC_5382 replaced by MAC_5826

//MAC_5393 replaced by MAC_5827

//MAC_5392 replaced by MAC_5827

//MAC_5391 replaced by MAC_5826

//MAC_5390 replaced by MAC_5827

//MAC_5389 replaced by MAC_5827

//MAC_5388 replaced by MAC_5826

//MAC_5399 replaced by MAC_5827

//MAC_5398 replaced by MAC_5827

//MAC_5397 replaced by MAC_5826

//MAC_5396 replaced by MAC_5827

//MAC_5395 replaced by MAC_5827

//MAC_5394 replaced by MAC_5826

//MAC_5405 replaced by MAC_5827

//MAC_5404 replaced by MAC_5827

//MAC_5403 replaced by MAC_5826

//MAC_5402 replaced by MAC_5827

//MAC_5401 replaced by MAC_5827

//MAC_5400 replaced by MAC_5826

//MAC_5411 replaced by MAC_5827

//MAC_5410 replaced by MAC_5827

//MAC_5409 replaced by MAC_5826

//MAC_5408 replaced by MAC_5827

//MAC_5407 replaced by MAC_5827

//MAC_5406 replaced by MAC_5826

//MAC_5417 replaced by MAC_5827

//MAC_5416 replaced by MAC_5827

//MAC_5415 replaced by MAC_5826

//MAC_5414 replaced by MAC_5827

//MAC_5413 replaced by MAC_5827

//MAC_5412 replaced by MAC_5826

//MAC_5423 replaced by MAC_5827

//MAC_5422 replaced by MAC_5827

//MAC_5421 replaced by MAC_5826

//MAC_5420 replaced by MAC_5827

//MAC_5419 replaced by MAC_5827

//MAC_5418 replaced by MAC_5826

//MAC_5429 replaced by MAC_5827

//MAC_5428 replaced by MAC_5827

//MAC_5427 replaced by MAC_5826

//MAC_5426 replaced by MAC_5827

//MAC_5425 replaced by MAC_5827

//MAC_5424 replaced by MAC_5826

//MAC_5435 replaced by MAC_5827

//MAC_5434 replaced by MAC_5827

//MAC_5433 replaced by MAC_5826

//MAC_5432 replaced by MAC_5827

//MAC_5431 replaced by MAC_5827

//MAC_5430 replaced by MAC_5826

//MAC_5441 replaced by MAC_5827

//MAC_5440 replaced by MAC_5827

//MAC_5439 replaced by MAC_5826

//MAC_5438 replaced by MAC_5827

//MAC_5437 replaced by MAC_5827

//MAC_5436 replaced by MAC_5826

//MAC_5447 replaced by MAC_5827

//MAC_5446 replaced by MAC_5827

//MAC_5445 replaced by MAC_5826

//MAC_5444 replaced by MAC_5827

//MAC_5443 replaced by MAC_5827

//MAC_5442 replaced by MAC_5826

//MAC_5453 replaced by MAC_5827

//MAC_5452 replaced by MAC_5827

//MAC_5451 replaced by MAC_5826

//MAC_5450 replaced by MAC_5827

//MAC_5449 replaced by MAC_5827

//MAC_5448 replaced by MAC_5826

//MAC_5459 replaced by MAC_5827

//MAC_5458 replaced by MAC_5827

//MAC_5457 replaced by MAC_5826

//MAC_5456 replaced by MAC_5827

//MAC_5455 replaced by MAC_5827

//MAC_5454 replaced by MAC_5826

//MAC_5465 replaced by MAC_5827

//MAC_5464 replaced by MAC_5827

//MAC_5463 replaced by MAC_5826

//MAC_5462 replaced by MAC_5827

//MAC_5461 replaced by MAC_5827

//MAC_5460 replaced by MAC_5826

//MAC_5471 replaced by MAC_5827

//MAC_5470 replaced by MAC_5827

//MAC_5469 replaced by MAC_5826

//MAC_5468 replaced by MAC_5827

//MAC_5467 replaced by MAC_5827

//MAC_5466 replaced by MAC_5826

//MAC_5477 replaced by MAC_5827

//MAC_5476 replaced by MAC_5827

//MAC_5475 replaced by MAC_5826

//MAC_5474 replaced by MAC_5827

//MAC_5473 replaced by MAC_5827

//MAC_5472 replaced by MAC_5826

//MAC_5483 replaced by MAC_5827

//MAC_5482 replaced by MAC_5827

//MAC_5481 replaced by MAC_5826

//MAC_5480 replaced by MAC_5827

//MAC_5479 replaced by MAC_5827

//MAC_5478 replaced by MAC_5826

//MAC_5489 replaced by MAC_5827

//MAC_5488 replaced by MAC_5827

//MAC_5487 replaced by MAC_5826

//MAC_5486 replaced by MAC_5827

//MAC_5485 replaced by MAC_5827

//MAC_5484 replaced by MAC_5826

//MAC_5495 replaced by MAC_5827

//MAC_5494 replaced by MAC_5827

//MAC_5493 replaced by MAC_5826

//MAC_5492 replaced by MAC_5827

//MAC_5491 replaced by MAC_5827

//MAC_5490 replaced by MAC_5826

//MAC_5501 replaced by MAC_5827

//MAC_5500 replaced by MAC_5827

//MAC_5499 replaced by MAC_5826

//MAC_5498 replaced by MAC_5827

//MAC_5497 replaced by MAC_5827

//MAC_5496 replaced by MAC_5826

//MAC_5507 replaced by MAC_5827

//MAC_5506 replaced by MAC_5827

//MAC_5505 replaced by MAC_5826

//MAC_5504 replaced by MAC_5827

//MAC_5503 replaced by MAC_5827

//MAC_5502 replaced by MAC_5826

//MAC_5513 replaced by MAC_5827

//MAC_5512 replaced by MAC_5827

//MAC_5511 replaced by MAC_5826

//MAC_5510 replaced by MAC_5827

//MAC_5509 replaced by MAC_5827

//MAC_5508 replaced by MAC_5826

//MAC_5519 replaced by MAC_5827

//MAC_5518 replaced by MAC_5827

//MAC_5517 replaced by MAC_5826

//MAC_5516 replaced by MAC_5827

//MAC_5515 replaced by MAC_5827

//MAC_5514 replaced by MAC_5826

//MAC_5525 replaced by MAC_5827

//MAC_5524 replaced by MAC_5827

//MAC_5523 replaced by MAC_5826

//MAC_5522 replaced by MAC_5827

//MAC_5521 replaced by MAC_5827

//MAC_5520 replaced by MAC_5826

//MAC_5531 replaced by MAC_5827

//MAC_5530 replaced by MAC_5827

//MAC_5529 replaced by MAC_5826

//MAC_5528 replaced by MAC_5827

//MAC_5527 replaced by MAC_5827

//MAC_5526 replaced by MAC_5826

//MAC_5537 replaced by MAC_5827

//MAC_5536 replaced by MAC_5827

//MAC_5535 replaced by MAC_5826

//MAC_5534 replaced by MAC_5827

//MAC_5533 replaced by MAC_5827

//MAC_5532 replaced by MAC_5826

//MAC_5543 replaced by MAC_5827

//MAC_5542 replaced by MAC_5827

//MAC_5541 replaced by MAC_5826

//MAC_5540 replaced by MAC_5827

//MAC_5539 replaced by MAC_5827

//MAC_5538 replaced by MAC_5826

//MAC_5549 replaced by MAC_5827

//MAC_5548 replaced by MAC_5827

//MAC_5547 replaced by MAC_5826

//MAC_5546 replaced by MAC_5827

//MAC_5545 replaced by MAC_5827

//MAC_5544 replaced by MAC_5826

//MAC_5555 replaced by MAC_5827

//MAC_5554 replaced by MAC_5827

//MAC_5553 replaced by MAC_5826

//MAC_5552 replaced by MAC_5827

//MAC_5551 replaced by MAC_5827

//MAC_5550 replaced by MAC_5826

//MAC_5561 replaced by MAC_5827

//MAC_5560 replaced by MAC_5827

//MAC_5559 replaced by MAC_5826

//MAC_5558 replaced by MAC_5827

//MAC_5557 replaced by MAC_5827

//MAC_5556 replaced by MAC_5826

//MAC_5567 replaced by MAC_5827

//MAC_5566 replaced by MAC_5827

//MAC_5565 replaced by MAC_5826

//MAC_5564 replaced by MAC_5827

//MAC_5563 replaced by MAC_5827

//MAC_5562 replaced by MAC_5826

//MAC_5573 replaced by MAC_5827

//MAC_5572 replaced by MAC_5827

//MAC_5571 replaced by MAC_5826

//MAC_5570 replaced by MAC_5827

//MAC_5569 replaced by MAC_5827

//MAC_5568 replaced by MAC_5826

//MAC_5579 replaced by MAC_5827

//MAC_5578 replaced by MAC_5827

//MAC_5577 replaced by MAC_5826

//MAC_5576 replaced by MAC_5827

//MAC_5575 replaced by MAC_5827

//MAC_5574 replaced by MAC_5826

//MAC_5585 replaced by MAC_5827

//MAC_5584 replaced by MAC_5827

//MAC_5583 replaced by MAC_5826

//MAC_5582 replaced by MAC_5827

//MAC_5581 replaced by MAC_5827

//MAC_5580 replaced by MAC_5826

//MAC_5591 replaced by MAC_5827

//MAC_5590 replaced by MAC_5827

//MAC_5589 replaced by MAC_5826

//MAC_5588 replaced by MAC_5827

//MAC_5587 replaced by MAC_5827

//MAC_5586 replaced by MAC_5826

//MAC_5597 replaced by MAC_5827

//MAC_5596 replaced by MAC_5827

//MAC_5595 replaced by MAC_5826

//MAC_5594 replaced by MAC_5827

//MAC_5593 replaced by MAC_5827

//MAC_5592 replaced by MAC_5826

//MAC_5603 replaced by MAC_5827

//MAC_5602 replaced by MAC_5827

//MAC_5601 replaced by MAC_5826

//MAC_5600 replaced by MAC_5827

//MAC_5599 replaced by MAC_5827

//MAC_5598 replaced by MAC_5826

//MAC_5609 replaced by MAC_5827

//MAC_5608 replaced by MAC_5827

//MAC_5607 replaced by MAC_5826

//MAC_5606 replaced by MAC_5827

//MAC_5605 replaced by MAC_5827

//MAC_5604 replaced by MAC_5826

//MAC_5615 replaced by MAC_5827

//MAC_5614 replaced by MAC_5827

//MAC_5613 replaced by MAC_5826

//MAC_5612 replaced by MAC_5827

//MAC_5611 replaced by MAC_5827

//MAC_5610 replaced by MAC_5826

//MAC_5621 replaced by MAC_5827

//MAC_5620 replaced by MAC_5827

//MAC_5619 replaced by MAC_5826

//MAC_5618 replaced by MAC_5827

//MAC_5617 replaced by MAC_5827

//MAC_5616 replaced by MAC_5826

//MAC_5627 replaced by MAC_5827

//MAC_5626 replaced by MAC_5827

//MAC_5625 replaced by MAC_5826

//MAC_5624 replaced by MAC_5827

//MAC_5623 replaced by MAC_5827

//MAC_5622 replaced by MAC_5826

//MAC_5633 replaced by MAC_5827

//MAC_5632 replaced by MAC_5827

//MAC_5631 replaced by MAC_5826

//MAC_5630 replaced by MAC_5827

//MAC_5629 replaced by MAC_5827

//MAC_5628 replaced by MAC_5826

//MAC_5639 replaced by MAC_5827

//MAC_5638 replaced by MAC_5827

//MAC_5637 replaced by MAC_5826

//MAC_5636 replaced by MAC_5827

//MAC_5635 replaced by MAC_5827

//MAC_5634 replaced by MAC_5826

//MAC_5645 replaced by MAC_5827

//MAC_5644 replaced by MAC_5827

//MAC_5643 replaced by MAC_5826

//MAC_5642 replaced by MAC_5827

//MAC_5641 replaced by MAC_5827

//MAC_5640 replaced by MAC_5826

//MAC_5651 replaced by MAC_5827

//MAC_5650 replaced by MAC_5827

//MAC_5649 replaced by MAC_5826

//MAC_5648 replaced by MAC_5827

//MAC_5647 replaced by MAC_5827

//MAC_5646 replaced by MAC_5826

//MAC_5657 replaced by MAC_5827

//MAC_5656 replaced by MAC_5827

//MAC_5655 replaced by MAC_5826

//MAC_5654 replaced by MAC_5827

//MAC_5653 replaced by MAC_5827

//MAC_5652 replaced by MAC_5826

//MAC_5663 replaced by MAC_5827

//MAC_5662 replaced by MAC_5827

//MAC_5661 replaced by MAC_5826

//MAC_5660 replaced by MAC_5827

//MAC_5659 replaced by MAC_5827

//MAC_5658 replaced by MAC_5826

//MAC_5669 replaced by MAC_5827

//MAC_5668 replaced by MAC_5827

//MAC_5667 replaced by MAC_5826

//MAC_5666 replaced by MAC_5827

//MAC_5665 replaced by MAC_5827

//MAC_5664 replaced by MAC_5826

//MAC_5675 replaced by MAC_5827

//MAC_5674 replaced by MAC_5827

//MAC_5673 replaced by MAC_5826

//MAC_5672 replaced by MAC_5827

//MAC_5671 replaced by MAC_5827

//MAC_5670 replaced by MAC_5826

//MAC_5681 replaced by MAC_5827

//MAC_5680 replaced by MAC_5827

//MAC_5679 replaced by MAC_5826

//MAC_5678 replaced by MAC_5827

//MAC_5677 replaced by MAC_5827

//MAC_5676 replaced by MAC_5826

//MAC_5687 replaced by MAC_5827

//MAC_5686 replaced by MAC_5827

//MAC_5685 replaced by MAC_5826

//MAC_5684 replaced by MAC_5827

//MAC_5683 replaced by MAC_5827

//MAC_5682 replaced by MAC_5826

//MAC_5693 replaced by MAC_5827

//MAC_5692 replaced by MAC_5827

//MAC_5691 replaced by MAC_5826

//MAC_5690 replaced by MAC_5827

//MAC_5689 replaced by MAC_5827

//MAC_5688 replaced by MAC_5826

//MAC_5699 replaced by MAC_5827

//MAC_5698 replaced by MAC_5827

//MAC_5697 replaced by MAC_5826

//MAC_5696 replaced by MAC_5827

//MAC_5695 replaced by MAC_5827

//MAC_5694 replaced by MAC_5826

//MAC_5705 replaced by MAC_5827

//MAC_5704 replaced by MAC_5827

//MAC_5703 replaced by MAC_5826

//MAC_5702 replaced by MAC_5827

//MAC_5701 replaced by MAC_5827

//MAC_5700 replaced by MAC_5826

//MAC_5711 replaced by MAC_5827

//MAC_5710 replaced by MAC_5827

//MAC_5709 replaced by MAC_5826

//MAC_5708 replaced by MAC_5827

//MAC_5707 replaced by MAC_5827

//MAC_5706 replaced by MAC_5826

//MAC_5717 replaced by MAC_5827

//MAC_5716 replaced by MAC_5827

//MAC_5715 replaced by MAC_5826

//MAC_5714 replaced by MAC_5827

//MAC_5713 replaced by MAC_5827

//MAC_5712 replaced by MAC_5826

//MAC_5723 replaced by MAC_5827

//MAC_5722 replaced by MAC_5827

//MAC_5721 replaced by MAC_5826

//MAC_5720 replaced by MAC_5827

//MAC_5719 replaced by MAC_5827

//MAC_5718 replaced by MAC_5826

//MAC_5729 replaced by MAC_5827

//MAC_5728 replaced by MAC_5827

//MAC_5727 replaced by MAC_5826

//MAC_5726 replaced by MAC_5827

//MAC_5725 replaced by MAC_5827

//MAC_5724 replaced by MAC_5826

//MAC_5735 replaced by MAC_5827

//MAC_5734 replaced by MAC_5827

//MAC_5733 replaced by MAC_5826

//MAC_5732 replaced by MAC_5827

//MAC_5731 replaced by MAC_5827

//MAC_5730 replaced by MAC_5826

//MAC_5741 replaced by MAC_5827

//MAC_5740 replaced by MAC_5827

//MAC_5739 replaced by MAC_5826

//MAC_5738 replaced by MAC_5827

//MAC_5737 replaced by MAC_5827

//MAC_5736 replaced by MAC_5826

//MAC_5747 replaced by MAC_5827

//MAC_5746 replaced by MAC_5827

//MAC_5745 replaced by MAC_5826

//MAC_5744 replaced by MAC_5827

//MAC_5743 replaced by MAC_5827

//MAC_5742 replaced by MAC_5826

//MAC_5753 replaced by MAC_5827

//MAC_5752 replaced by MAC_5827

//MAC_5751 replaced by MAC_5826

//MAC_5750 replaced by MAC_5827

//MAC_5749 replaced by MAC_5827

//MAC_5748 replaced by MAC_5826

//MAC_5759 replaced by MAC_5827

//MAC_5758 replaced by MAC_5827

//MAC_5757 replaced by MAC_5826

//MAC_5756 replaced by MAC_5827

//MAC_5755 replaced by MAC_5827

//MAC_5754 replaced by MAC_5826

//MAC_5765 replaced by MAC_5827

//MAC_5764 replaced by MAC_5827

//MAC_5763 replaced by MAC_5826

//MAC_5762 replaced by MAC_5827

//MAC_5761 replaced by MAC_5827

//MAC_5760 replaced by MAC_5826

//MAC_5771 replaced by MAC_5827

//MAC_5770 replaced by MAC_5827

//MAC_5769 replaced by MAC_5826

//MAC_5768 replaced by MAC_5827

//MAC_5767 replaced by MAC_5827

//MAC_5766 replaced by MAC_5826

//MAC_5777 replaced by MAC_5827

//MAC_5776 replaced by MAC_5827

//MAC_5775 replaced by MAC_5826

//MAC_5774 replaced by MAC_5827

//MAC_5773 replaced by MAC_5827

//MAC_5772 replaced by MAC_5826

//MAC_5783 replaced by MAC_5827

//MAC_5782 replaced by MAC_5827

//MAC_5781 replaced by MAC_5826

//MAC_5780 replaced by MAC_5827

//MAC_5779 replaced by MAC_5827

//MAC_5778 replaced by MAC_5826

//MAC_5789 replaced by MAC_5827

//MAC_5788 replaced by MAC_5827

//MAC_5787 replaced by MAC_5826

//MAC_5786 replaced by MAC_5827

//MAC_5785 replaced by MAC_5827

//MAC_5784 replaced by MAC_5826

//MAC_5795 replaced by MAC_5827

//MAC_5794 replaced by MAC_5827

//MAC_5793 replaced by MAC_5826

//MAC_5792 replaced by MAC_5827

//MAC_5791 replaced by MAC_5827

//MAC_5790 replaced by MAC_5826

//MAC_5801 replaced by MAC_5827

//MAC_5800 replaced by MAC_5827

//MAC_5799 replaced by MAC_5826

//MAC_5798 replaced by MAC_5827

//MAC_5797 replaced by MAC_5827

//MAC_5796 replaced by MAC_5826

//MAC_5807 replaced by MAC_5827

//MAC_5806 replaced by MAC_5827

//MAC_5805 replaced by MAC_5826

//MAC_5804 replaced by MAC_5827

//MAC_5803 replaced by MAC_5827

//MAC_5802 replaced by MAC_5826

//MAC_5813 replaced by MAC_5827

//MAC_5812 replaced by MAC_5827

//MAC_5811 replaced by MAC_5826

//MAC_5810 replaced by MAC_5827

//MAC_5809 replaced by MAC_5827

//MAC_5808 replaced by MAC_5826

//MAC_5819 replaced by MAC_5827

//MAC_5818 replaced by MAC_5827

//MAC_5817 replaced by MAC_5826

//MAC_5816 replaced by MAC_5827

//MAC_5815 replaced by MAC_5827

//MAC_5814 replaced by MAC_5826

//MAC_5825 replaced by MAC_5827

//MAC_5824 replaced by MAC_5827

//MAC_5823 replaced by MAC_5826

//MAC_5822 replaced by MAC_5827

//MAC_5821 replaced by MAC_5827

//MAC_5820 replaced by MAC_5826

//MAC_5831 replaced by MAC_5827

//MAC_5830 replaced by MAC_5827

//MAC_5829 replaced by MAC_5826

//MAC_5828 replaced by MAC_5827

module MAC_5827 (
  input      [25:0]   io_a,
  input      [29:0]   io_acin,
  output     [29:0]   io_acout,
  input      [16:0]   io_b,
  input      [16:0]   io_c,
  input               io_ce,
  input      [47:0]   io_pcin,
  output     [42:0]   io_p,
  output     [47:0]   io_pcout,
  input               clk
);

  wire       [29:0]   DSP_A;
  wire       [17:0]   DSP_B;
  wire       [47:0]   DSP_C;
  wire       [8:0]    DSP_OPMODE;
  wire       [29:0]   DSP_ACOUT;
  wire       [47:0]   DSP_P;
  wire       [47:0]   DSP_PCOUT;
  wire       [26:0]   _zz_A;
  wire       [0:0]    _zz_A_1;
  wire       [0:0]    _zz_B;
  wire       [17:0]   _zz_C;
  wire       [0:0]    _zz_C_1;
  wire       [47:0]   _zz_io_p;

  assign _zz_A = {_zz_A_1,io_a};
  assign _zz_A_1 = 1'b0;
  assign _zz_B = 1'b0;
  assign _zz_C = {_zz_C_1,io_c};
  assign _zz_C_1 = 1'b0;
  assign _zz_io_p = DSP_P;
  DSP48E2 #(
    .A_INPUT("CASCADE"),
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AMULTSEL("A"),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .AUTORESET_PRIORITY("RESET"),
    .B_INPUT ("DIRECT"),
    .BCASCREG(1),
    .BMULTSEL("B"),
    .BREG(1),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'h0),
    .IS_OPMODE_INVERTED(9'h0),
    .IS_RSTA_INVERTED(1'b0),
    .IS_RSTALLCARRYIN_INVERTED(1'b0),
    .IS_RSTALUMODE_INVERTED(1'b0),
    .IS_RSTB_INVERTED(1'b0),
    .IS_RSTC_INVERTED(1'b0),
    .IS_RSTCTRL_INVERTED(1'b0),
    .IS_RSTD_INVERTED(1'b0),
    .IS_RSTINMODE_INVERTED(1'b0),
    .IS_RSTM_INVERTED(1'b0),
    .IS_RSTP_INVERTED(1'b0),
    .MASK(48'h0),
    .MREG(1),
    .OPMODEREG(1),
    .PATTERN(48'h0),
    .PREADDINSEL("A"),
    .PREG(1),
    .RND(48'h0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48"),
    .USE_WIDEXOR("FALSE"),
    .XORSIMD("XOR24_48_96")
  ) DSP (
    .A             (DSP_A[29:0]    ), //i
    .ACIN          (io_acin[29:0]  ), //i
    .ACOUT         (DSP_ACOUT[29:0]), //o
    .B             (DSP_B[17:0]    ), //i
    .C             (DSP_C[47:0]    ), //i
    .CLK           (clk            ), //i
    .OPMODE        (DSP_OPMODE[8:0]), //i
    .P             (DSP_P[47:0]    ), //o
    .PCIN          (io_pcin[47:0]  ), //i
    .PCOUT         (DSP_PCOUT[47:0]), //o
    .ALUMODE       (4'b0000        ), //i
    .BCIN          (18'h0          ), //i
    .CARRYCASCIN   (1'b0           ), //i
    .CARRYIN       (1'b0           ), //i
    .CARRYINSEL    (3'b000         ), //i
    .CEA1          (1'b0           ), //i
    .CEA2          (1'b1           ), //i
    .CEAD          (1'b0           ), //i
    .CEALUMODE     (1'b0           ), //i
    .CEB1          (1'b0           ), //i
    .CEB2          (1'b1           ), //i
    .CEC           (1'b1           ), //i
    .CECARRYIN     (1'b0           ), //i
    .CECTRL        (1'b1           ), //i
    .CED           (1'b0           ), //i
    .CEINMODE      (1'b0           ), //i
    .CEM           (1'b1           ), //i
    .CEP           (1'b1           ), //i
    .D             (27'h0          ), //i
    .INMODE        (5'h0           ), //i
    .MULTSIGNIN    (1'b0           ), //i
    .RSTA          (1'b0           ), //i
    .RSTALLCARRYIN (1'b0           ), //i
    .RSTALUMODE    (1'b0           ), //i
    .RSTB          (1'b0           ), //i
    .RSTC          (1'b0           ), //i
    .RSTCTRL       (1'b0           ), //i
    .RSTD          (1'b0           ), //i
    .RSTINMODE     (1'b0           ), //i
    .RSTM          (1'b0           ), //i
    .RSTP          (1'b0           )  //i
  );
  assign DSP_A = {{3{_zz_A[26]}}, _zz_A};
  assign io_acout = DSP_ACOUT;
  assign DSP_B = {_zz_B,io_b};
  assign DSP_C = {{30{_zz_C[17]}}, _zz_C};
  assign DSP_OPMODE = {{io_ce,io_ce},7'h55};
  assign io_p = _zz_io_p[42:0];
  assign io_pcout = DSP_PCOUT;

endmodule

module MAC_5826 (
  input      [25:0]   io_a,
  input      [29:0]   io_acin,
  output     [29:0]   io_acout,
  input      [16:0]   io_b,
  input      [16:0]   io_c,
  input               io_ce,
  input      [47:0]   io_pcin,
  output     [42:0]   io_p,
  output     [47:0]   io_pcout,
  input               clk
);

  wire       [29:0]   DSP_A;
  wire       [17:0]   DSP_B;
  wire       [47:0]   DSP_C;
  wire       [8:0]    DSP_OPMODE;
  wire       [29:0]   DSP_ACOUT;
  wire       [47:0]   DSP_P;
  wire       [47:0]   DSP_PCOUT;
  wire       [26:0]   _zz_A;
  wire       [0:0]    _zz_A_1;
  wire       [0:0]    _zz_B;
  wire       [17:0]   _zz_C;
  wire       [0:0]    _zz_C_1;
  wire       [47:0]   _zz_io_p;

  assign _zz_A = {_zz_A_1,io_a};
  assign _zz_A_1 = 1'b0;
  assign _zz_B = 1'b0;
  assign _zz_C = {_zz_C_1,io_c};
  assign _zz_C_1 = 1'b0;
  assign _zz_io_p = DSP_P;
  DSP48E2 #(
    .A_INPUT("DIRECT"),
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AMULTSEL("A"),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .AUTORESET_PRIORITY("RESET"),
    .B_INPUT ("DIRECT"),
    .BCASCREG(1),
    .BMULTSEL("B"),
    .BREG(1),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'h0),
    .IS_OPMODE_INVERTED(9'h0),
    .IS_RSTA_INVERTED(1'b0),
    .IS_RSTALLCARRYIN_INVERTED(1'b0),
    .IS_RSTALUMODE_INVERTED(1'b0),
    .IS_RSTB_INVERTED(1'b0),
    .IS_RSTC_INVERTED(1'b0),
    .IS_RSTCTRL_INVERTED(1'b0),
    .IS_RSTD_INVERTED(1'b0),
    .IS_RSTINMODE_INVERTED(1'b0),
    .IS_RSTM_INVERTED(1'b0),
    .IS_RSTP_INVERTED(1'b0),
    .MASK(48'h0),
    .MREG(1),
    .OPMODEREG(1),
    .PATTERN(48'h0),
    .PREADDINSEL("A"),
    .PREG(1),
    .RND(48'h0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48"),
    .USE_WIDEXOR("FALSE"),
    .XORSIMD("XOR24_48_96")
  ) DSP (
    .A             (DSP_A[29:0]    ), //i
    .ACIN          (io_acin[29:0]  ), //i
    .ACOUT         (DSP_ACOUT[29:0]), //o
    .B             (DSP_B[17:0]    ), //i
    .C             (DSP_C[47:0]    ), //i
    .CLK           (clk            ), //i
    .OPMODE        (DSP_OPMODE[8:0]), //i
    .P             (DSP_P[47:0]    ), //o
    .PCIN          (io_pcin[47:0]  ), //i
    .PCOUT         (DSP_PCOUT[47:0]), //o
    .ALUMODE       (4'b0000        ), //i
    .BCIN          (18'h0          ), //i
    .CARRYCASCIN   (1'b0           ), //i
    .CARRYIN       (1'b0           ), //i
    .CARRYINSEL    (3'b000         ), //i
    .CEA1          (1'b0           ), //i
    .CEA2          (1'b1           ), //i
    .CEAD          (1'b0           ), //i
    .CEALUMODE     (1'b0           ), //i
    .CEB1          (1'b0           ), //i
    .CEB2          (1'b1           ), //i
    .CEC           (1'b1           ), //i
    .CECARRYIN     (1'b0           ), //i
    .CECTRL        (1'b1           ), //i
    .CED           (1'b0           ), //i
    .CEINMODE      (1'b0           ), //i
    .CEM           (1'b1           ), //i
    .CEP           (1'b1           ), //i
    .D             (27'h0          ), //i
    .INMODE        (5'h0           ), //i
    .MULTSIGNIN    (1'b0           ), //i
    .RSTA          (1'b0           ), //i
    .RSTALLCARRYIN (1'b0           ), //i
    .RSTALUMODE    (1'b0           ), //i
    .RSTB          (1'b0           ), //i
    .RSTC          (1'b0           ), //i
    .RSTCTRL       (1'b0           ), //i
    .RSTD          (1'b0           ), //i
    .RSTINMODE     (1'b0           ), //i
    .RSTM          (1'b0           ), //i
    .RSTP          (1'b0           )  //i
  );
  assign DSP_A = {{3{_zz_A[26]}}, _zz_A};
  assign io_acout = DSP_ACOUT;
  assign DSP_B = {_zz_B,io_b};
  assign DSP_C = {{30{_zz_C[17]}}, _zz_C};
  assign DSP_OPMODE = {{io_ce,io_ce},7'h05};
  assign io_p = _zz_io_p[42:0];
  assign io_pcout = DSP_PCOUT;

endmodule
