// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : PippengerU250
// Git hash  : d6da632995922518897eb20accafd73e16698ecf

`timescale 1ns/1ps

module PippengerU250 (
  output              dataBus_awvalid,
  input               dataBus_awready,
  output     [63:0]   dataBus_awaddr,
  output     [7:0]    dataBus_awlen,
  output              dataBus_wvalid,
  input               dataBus_wready,
  output     [511:0]  dataBus_wdata,
  output              dataBus_wlast,
  input               dataBus_bvalid,
  output              dataBus_bready,
  output              dataBus_arvalid,
  input               dataBus_arready,
  output     [63:0]   dataBus_araddr,
  output     [7:0]    dataBus_arlen,
  input               dataBus_rvalid,
  output              dataBus_rready,
  input      [511:0]  dataBus_rdata,
  input               dataBus_rlast,
  input               s_axi_control_awvalid,
  output              s_axi_control_awready,
  input      [5:0]    s_axi_control_awaddr,
  input      [2:0]    s_axi_control_awprot,
  input               s_axi_control_wvalid,
  output              s_axi_control_wready,
  input      [31:0]   s_axi_control_wdata,
  input      [3:0]    s_axi_control_wstrb,
  output              s_axi_control_bvalid,
  input               s_axi_control_bready,
  output     [1:0]    s_axi_control_bresp,
  input               s_axi_control_arvalid,
  output reg          s_axi_control_arready,
  input      [5:0]    s_axi_control_araddr,
  input      [2:0]    s_axi_control_arprot,
  output              s_axi_control_rvalid,
  input               s_axi_control_rready,
  output     [31:0]   s_axi_control_rdata,
  output     [1:0]    s_axi_control_rresp,
  input               clk,
  input               resetn
);

  wire       [376:0]  pippenger_1_io_dataIn_payload_fragment_P_X;
  wire       [376:0]  pippenger_1_io_dataIn_payload_fragment_P_Y;
  wire       [376:0]  pippenger_1_io_dataIn_payload_fragment_P_T;
  wire       [252:0]  pippenger_1_io_dataIn_payload_fragment_K;
  wire                dataBusReadArea_inputDMA_io_streamBus_ready;
  wire                pippenger_1_io_dataIn_ready;
  wire                pippenger_1_io_dataOut_valid;
  wire       [376:0]  pippenger_1_io_dataOut_payload_X;
  wire       [376:0]  pippenger_1_io_dataOut_payload_Y;
  wire       [376:0]  pippenger_1_io_dataOut_payload_Z;
  wire       [376:0]  pippenger_1_io_dataOut_payload_T;
  wire                dataBusReadArea_inputDMA_io_axi4Bus_ar_valid;
  wire       [63:0]   dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_addr;
  wire       [7:0]    dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_len;
  wire                dataBusReadArea_inputDMA_io_axi4Bus_r_ready;
  wire                dataBusReadArea_inputDMA_io_streamBus_valid;
  wire       [511:0]  dataBusReadArea_inputDMA_io_streamBus_payload;
  wire                dataBusReadArea_inputDMA_io_done;
  wire       [27:0]   _zz_pageNum;
  wire       [27:0]   _zz_pageNum_1;
  wire       [26:0]   _zz_pageNum_2;
  wire       [26:0]   _zz_pageNum_3;
  wire       [1:0]    _zz_dataBusReadArea_inputCnt_valueNext;
  wire       [0:0]    _zz_dataBusReadArea_inputCnt_valueNext_1;
  wire       [31:0]   _zz_dataBusReadArea_lastCnt_valueNext;
  wire       [0:0]    _zz_dataBusReadArea_lastCnt_valueNext_1;
  wire       [1:0]    _zz_dataBusWriteArea_outputCnt_valueNext;
  wire       [0:0]    _zz_dataBusWriteArea_outputCnt_valueNext_1;
  wire       [376:0]  _zz_dataBus_wdata;
  wire       [31:0]   _zz_startReadAddress;
  wire       [31:0]   _zz_startReadAddress_1;
  wire       [31:0]   _zz_startReadAddress_2;
  wire       [31:0]   _zz_startReadAddress_3;
  wire       [31:0]   _zz_startWriteAddress;
  wire       [31:0]   _zz_startWriteAddress_1;
  wire       [31:0]   _zz_startWriteAddress_2;
  wire       [31:0]   _zz_startWriteAddress_3;
  reg                 startRise;
  reg                 readStart;
  reg                 writeStart;
  reg        [25:0]   num;
  reg        [27:0]   pageNum;
  reg        [63:0]   startReadAddress;
  reg        [63:0]   startWriteAddress;
  wire                slaveFactory_readErrorFlag;
  wire                slaveFactory_writeErrorFlag;
  wire                slaveFactory_readHaltRequest;
  wire                slaveFactory_writeHaltRequest;
  wire                slaveFactory_writeJoinEvent_valid;
  wire                slaveFactory_writeJoinEvent_ready;
  wire                slaveFactory_writeJoinEvent_fire;
  reg        [1:0]    slaveFactory_writeRsp_resp;
  wire                slaveFactory_writeJoinEvent_translated_valid;
  wire                slaveFactory_writeJoinEvent_translated_ready;
  wire       [1:0]    slaveFactory_writeJoinEvent_translated_payload_resp;
  wire                _zz_slaveFactory_writeJoinEvent_translated_ready;
  reg                 _zz_slaveFactory_writeJoinEvent_translated_ready_1;
  wire                _zz_s_axi_control_bvalid;
  reg                 _zz_s_axi_control_bvalid_1;
  reg        [1:0]    _zz_s_axi_control_bresp;
  wire                when_Stream_l368;
  wire                slaveFactory_readDataStage_valid;
  wire                slaveFactory_readDataStage_ready;
  wire       [5:0]    slaveFactory_readDataStage_payload_addr;
  wire       [2:0]    slaveFactory_readDataStage_payload_prot;
  reg                 io_s_axi_control_ar_rValid;
  reg        [5:0]    io_s_axi_control_ar_rData_addr;
  reg        [2:0]    io_s_axi_control_ar_rData_prot;
  wire                when_Stream_l368_1;
  reg        [31:0]   slaveFactory_readRsp_data;
  reg        [1:0]    slaveFactory_readRsp_resp;
  wire                _zz_s_axi_control_rvalid;
  wire       [5:0]    slaveFactory_readAddressMasked;
  wire       [5:0]    slaveFactory_writeAddressMasked;
  wire                slaveFactory_writeOccur;
  wire                slaveFactory_readOccur;
  wire       [63:0]   _zz_slaveFactory_readRsp_data;
  wire       [63:0]   _zz_slaveFactory_readRsp_data_1;
  reg                 dataBusReadArea_inputCnt_willIncrement;
  wire                dataBusReadArea_inputCnt_willClear;
  reg        [1:0]    dataBusReadArea_inputCnt_valueNext;
  reg        [1:0]    dataBusReadArea_inputCnt_value;
  reg                 dataBusReadArea_inputCnt_willOverflowIfInc;
  wire                dataBusReadArea_inputCnt_willOverflow;
  reg                 dataBusReadArea_inputValid;
  reg        [511:0]  dataBusReadArea_inputData_0;
  reg        [511:0]  dataBusReadArea_inputData_1;
  reg        [511:0]  dataBusReadArea_inputData_2;
  wire       [383:0]  dataBusReadArea_outputData_0;
  wire       [383:0]  dataBusReadArea_outputData_1;
  wire       [383:0]  dataBusReadArea_outputData_2;
  wire       [383:0]  dataBusReadArea_outputData_3;
  wire       [1535:0] _zz_dataBusReadArea_outputData_0;
  reg                 dataBusReadArea_lastCnt_willIncrement;
  reg                 dataBusReadArea_lastCnt_willClear;
  reg        [31:0]   dataBusReadArea_lastCnt_valueNext;
  reg        [31:0]   dataBusReadArea_lastCnt_value;
  reg                 dataBusReadArea_lastCnt_willOverflowIfInc;
  wire                dataBusReadArea_lastCnt_willOverflow;
  wire                toplevel_pippenger_1_io_dataIn_fire;
  reg                 _zz_1;
  reg                 _zz_io_dataIn_payload_last;
  wire                toplevel_dataBusReadArea_inputDMA_io_streamBus_fire;
  reg                 dataBusWriteArea_outputCnt_willIncrement;
  wire                dataBusWriteArea_outputCnt_willClear;
  reg        [1:0]    dataBusWriteArea_outputCnt_valueNext;
  reg        [1:0]    dataBusWriteArea_outputCnt_value;
  reg                 dataBusWriteArea_outputCnt_willOverflowIfInc;
  wire                dataBusWriteArea_outputCnt_willOverflow;
  reg                 dataBusWriteArea_dataOutputValid;
  reg        [376:0]  dataBusWriteArea_dataReg_0;
  reg        [376:0]  dataBusWriteArea_dataReg_1;
  reg        [376:0]  dataBusWriteArea_dataReg_2;
  reg        [376:0]  dataBusWriteArea_dataReg_3;
  reg                 dataBusWriteArea_addressOutputValid;
  wire                io_dataBus_w_fire;
  wire                when_AxiLite4SlaveFactory_l68;
  wire                when_AxiLite4SlaveFactory_l68_1;
  wire                when_AxiLite4SlaveFactory_l68_2;
  wire                when_AxiLite4SlaveFactory_l68_3;
  wire                when_AxiLite4SlaveFactory_l86;
  wire                when_AxiLite4SlaveFactory_l86_1;
  wire                when_AxiLite4SlaveFactory_l86_2;
  wire                when_AxiLite4SlaveFactory_l86_3;

  assign _zz_pageNum = (_zz_pageNum_1 + {1'b0,_zz_pageNum_3});
  assign _zz_pageNum_2 = {1'b0,num};
  assign _zz_pageNum_1 = {1'd0, _zz_pageNum_2};
  assign _zz_pageNum_3 = ({1'd0,num} <<< 1);
  assign _zz_dataBusReadArea_inputCnt_valueNext_1 = dataBusReadArea_inputCnt_willIncrement;
  assign _zz_dataBusReadArea_inputCnt_valueNext = {1'd0, _zz_dataBusReadArea_inputCnt_valueNext_1};
  assign _zz_dataBusReadArea_lastCnt_valueNext_1 = dataBusReadArea_lastCnt_willIncrement;
  assign _zz_dataBusReadArea_lastCnt_valueNext = {31'd0, _zz_dataBusReadArea_lastCnt_valueNext_1};
  assign _zz_dataBusWriteArea_outputCnt_valueNext_1 = dataBusWriteArea_outputCnt_willIncrement;
  assign _zz_dataBusWriteArea_outputCnt_valueNext = {1'd0, _zz_dataBusWriteArea_outputCnt_valueNext_1};
  assign _zz_dataBus_wdata = dataBusWriteArea_dataReg_0;
  assign _zz_startReadAddress_1 = s_axi_control_wdata[31 : 0];
  assign _zz_startReadAddress = _zz_startReadAddress_1;
  assign _zz_startReadAddress_3 = s_axi_control_wdata[31 : 0];
  assign _zz_startReadAddress_2 = _zz_startReadAddress_3;
  assign _zz_startWriteAddress_1 = s_axi_control_wdata[31 : 0];
  assign _zz_startWriteAddress = _zz_startWriteAddress_1;
  assign _zz_startWriteAddress_3 = s_axi_control_wdata[31 : 0];
  assign _zz_startWriteAddress_2 = _zz_startWriteAddress_3;
  PippengerWithPAdd pippenger_1 (
    .io_dataIn_valid                (dataBusReadArea_inputValid                                                                          ), //i
    .io_dataIn_ready                (pippenger_1_io_dataIn_ready                                                                         ), //o
    .io_dataIn_payload_last         (_zz_io_dataIn_payload_last                                                                          ), //i
    .io_dataIn_payload_fragment_P_X (pippenger_1_io_dataIn_payload_fragment_P_X[376:0]                                                   ), //i
    .io_dataIn_payload_fragment_P_Y (pippenger_1_io_dataIn_payload_fragment_P_Y[376:0]                                                   ), //i
    .io_dataIn_payload_fragment_P_Z (377'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001), //i
    .io_dataIn_payload_fragment_P_T (pippenger_1_io_dataIn_payload_fragment_P_T[376:0]                                                   ), //i
    .io_dataIn_payload_fragment_K   (pippenger_1_io_dataIn_payload_fragment_K[252:0]                                                     ), //i
    .io_dataOut_valid               (pippenger_1_io_dataOut_valid                                                                        ), //o
    .io_dataOut_ready               (1'b1                                                                                                ), //i
    .io_dataOut_payload_X           (pippenger_1_io_dataOut_payload_X[376:0]                                                             ), //o
    .io_dataOut_payload_Y           (pippenger_1_io_dataOut_payload_Y[376:0]                                                             ), //o
    .io_dataOut_payload_Z           (pippenger_1_io_dataOut_payload_Z[376:0]                                                             ), //o
    .io_dataOut_payload_T           (pippenger_1_io_dataOut_payload_T[376:0]                                                             ), //o
    .clk                            (clk                                                                                                 ), //i
    .resetn                         (resetn                                                                                              )  //i
  );
  Axi4PageRDMA dataBusReadArea_inputDMA (
    .io_axi4Bus_ar_valid        (dataBusReadArea_inputDMA_io_axi4Bus_ar_valid             ), //o
    .io_axi4Bus_ar_ready        (dataBus_arready                                          ), //i
    .io_axi4Bus_ar_payload_addr (dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_addr[63:0]), //o
    .io_axi4Bus_ar_payload_len  (dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_len[7:0]  ), //o
    .io_axi4Bus_r_valid         (dataBus_rvalid                                           ), //i
    .io_axi4Bus_r_ready         (dataBusReadArea_inputDMA_io_axi4Bus_r_ready              ), //o
    .io_axi4Bus_r_payload_data  (dataBus_rdata[511:0]                                     ), //i
    .io_axi4Bus_r_payload_last  (dataBus_rlast                                            ), //i
    .io_streamBus_valid         (dataBusReadArea_inputDMA_io_streamBus_valid              ), //o
    .io_streamBus_ready         (dataBusReadArea_inputDMA_io_streamBus_ready              ), //i
    .io_streamBus_payload       (dataBusReadArea_inputDMA_io_streamBus_payload[511:0]     ), //o
    .io_work                    (readStart                                                ), //i
    .io_address                 (startReadAddress[63:0]                                   ), //i
    .io_pageNum                 (pageNum[27:0]                                            ), //i
    .io_done                    (dataBusReadArea_inputDMA_io_done                         ), //o
    .clk                        (clk                                                      ), //i
    .resetn                     (resetn                                                   )  //i
  );
  always @(*) begin
    startRise = 1'b0;
    case(slaveFactory_writeAddressMasked)
      6'h10 : begin
        if(slaveFactory_writeOccur) begin
          startRise = s_axi_control_wdata[0];
        end
      end
      default : begin
      end
    endcase
  end

  assign slaveFactory_readErrorFlag = 1'b0;
  assign slaveFactory_writeErrorFlag = 1'b0;
  assign slaveFactory_readHaltRequest = 1'b0;
  assign slaveFactory_writeHaltRequest = 1'b0;
  assign slaveFactory_writeJoinEvent_fire = (slaveFactory_writeJoinEvent_valid && slaveFactory_writeJoinEvent_ready);
  assign slaveFactory_writeJoinEvent_valid = (s_axi_control_awvalid && s_axi_control_wvalid);
  assign s_axi_control_awready = slaveFactory_writeJoinEvent_fire;
  assign s_axi_control_wready = slaveFactory_writeJoinEvent_fire;
  assign slaveFactory_writeJoinEvent_translated_valid = slaveFactory_writeJoinEvent_valid;
  assign slaveFactory_writeJoinEvent_ready = slaveFactory_writeJoinEvent_translated_ready;
  assign slaveFactory_writeJoinEvent_translated_payload_resp = slaveFactory_writeRsp_resp;
  assign _zz_slaveFactory_writeJoinEvent_translated_ready = (! slaveFactory_writeHaltRequest);
  assign slaveFactory_writeJoinEvent_translated_ready = (_zz_slaveFactory_writeJoinEvent_translated_ready_1 && _zz_slaveFactory_writeJoinEvent_translated_ready);
  always @(*) begin
    _zz_slaveFactory_writeJoinEvent_translated_ready_1 = s_axi_control_bready;
    if(when_Stream_l368) begin
      _zz_slaveFactory_writeJoinEvent_translated_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l368 = (! _zz_s_axi_control_bvalid);
  assign _zz_s_axi_control_bvalid = _zz_s_axi_control_bvalid_1;
  assign s_axi_control_bvalid = _zz_s_axi_control_bvalid;
  assign s_axi_control_bresp = _zz_s_axi_control_bresp;
  always @(*) begin
    s_axi_control_arready = slaveFactory_readDataStage_ready;
    if(when_Stream_l368_1) begin
      s_axi_control_arready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! slaveFactory_readDataStage_valid);
  assign slaveFactory_readDataStage_valid = io_s_axi_control_ar_rValid;
  assign slaveFactory_readDataStage_payload_addr = io_s_axi_control_ar_rData_addr;
  assign slaveFactory_readDataStage_payload_prot = io_s_axi_control_ar_rData_prot;
  assign _zz_s_axi_control_rvalid = (! slaveFactory_readHaltRequest);
  assign slaveFactory_readDataStage_ready = (s_axi_control_rready && _zz_s_axi_control_rvalid);
  assign s_axi_control_rvalid = (slaveFactory_readDataStage_valid && _zz_s_axi_control_rvalid);
  assign s_axi_control_rdata = slaveFactory_readRsp_data;
  assign s_axi_control_rresp = slaveFactory_readRsp_resp;
  always @(*) begin
    if(slaveFactory_writeErrorFlag) begin
      slaveFactory_writeRsp_resp = 2'b10;
    end else begin
      slaveFactory_writeRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    if(slaveFactory_readErrorFlag) begin
      slaveFactory_readRsp_resp = 2'b10;
    end else begin
      slaveFactory_readRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    slaveFactory_readRsp_data = 32'h0;
    case(slaveFactory_readAddressMasked)
      6'h10 : begin
        slaveFactory_readRsp_data[0 : 0] = (readStart || writeStart);
      end
      6'h18 : begin
        slaveFactory_readRsp_data[31 : 0] = {num,6'h3f};
      end
      default : begin
      end
    endcase
    if(when_AxiLite4SlaveFactory_l86) begin
      slaveFactory_readRsp_data[31 : 0] = _zz_slaveFactory_readRsp_data[31 : 0];
    end
    if(when_AxiLite4SlaveFactory_l86_1) begin
      slaveFactory_readRsp_data[31 : 0] = _zz_slaveFactory_readRsp_data[63 : 32];
    end
    if(when_AxiLite4SlaveFactory_l86_2) begin
      slaveFactory_readRsp_data[31 : 0] = _zz_slaveFactory_readRsp_data_1[31 : 0];
    end
    if(when_AxiLite4SlaveFactory_l86_3) begin
      slaveFactory_readRsp_data[31 : 0] = _zz_slaveFactory_readRsp_data_1[63 : 32];
    end
  end

  assign slaveFactory_readAddressMasked = (slaveFactory_readDataStage_payload_addr & (~ 6'h03));
  assign slaveFactory_writeAddressMasked = (s_axi_control_awaddr & (~ 6'h03));
  assign slaveFactory_writeOccur = (slaveFactory_writeJoinEvent_valid && slaveFactory_writeJoinEvent_ready);
  assign slaveFactory_readOccur = (s_axi_control_rvalid && s_axi_control_rready);
  assign _zz_slaveFactory_readRsp_data = startReadAddress;
  assign _zz_slaveFactory_readRsp_data_1 = startWriteAddress;
  assign dataBus_arvalid = dataBusReadArea_inputDMA_io_axi4Bus_ar_valid;
  assign dataBus_araddr = dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_addr;
  assign dataBus_arlen = dataBusReadArea_inputDMA_io_axi4Bus_ar_payload_len;
  assign dataBus_rready = dataBusReadArea_inputDMA_io_axi4Bus_r_ready;
  always @(*) begin
    dataBusReadArea_inputCnt_willIncrement = 1'b0;
    if(toplevel_dataBusReadArea_inputDMA_io_streamBus_fire) begin
      dataBusReadArea_inputCnt_willIncrement = 1'b1;
    end
  end

  assign dataBusReadArea_inputCnt_willClear = 1'b0;
  assign dataBusReadArea_inputCnt_willOverflow = (dataBusReadArea_inputCnt_willOverflowIfInc && dataBusReadArea_inputCnt_willIncrement);
  always @(*) begin
    if(dataBusReadArea_inputCnt_willOverflow) begin
      dataBusReadArea_inputCnt_valueNext = 2'b00;
    end else begin
      dataBusReadArea_inputCnt_valueNext = (dataBusReadArea_inputCnt_value + _zz_dataBusReadArea_inputCnt_valueNext);
    end
    if(dataBusReadArea_inputCnt_willClear) begin
      dataBusReadArea_inputCnt_valueNext = 2'b00;
    end
  end

  assign _zz_dataBusReadArea_outputData_0 = {dataBusReadArea_inputData_2,{dataBusReadArea_inputData_1,dataBusReadArea_inputData_0}};
  assign dataBusReadArea_outputData_0 = _zz_dataBusReadArea_outputData_0[383 : 0];
  assign dataBusReadArea_outputData_1 = _zz_dataBusReadArea_outputData_0[767 : 384];
  assign dataBusReadArea_outputData_2 = _zz_dataBusReadArea_outputData_0[1151 : 768];
  assign dataBusReadArea_outputData_3 = _zz_dataBusReadArea_outputData_0[1535 : 1152];
  always @(*) begin
    dataBusReadArea_lastCnt_willIncrement = 1'b0;
    if(toplevel_pippenger_1_io_dataIn_fire) begin
      dataBusReadArea_lastCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    dataBusReadArea_lastCnt_willClear = 1'b0;
    if(toplevel_pippenger_1_io_dataIn_fire) begin
      if(_zz_1) begin
        dataBusReadArea_lastCnt_willClear = 1'b1;
      end
    end
  end

  assign dataBusReadArea_lastCnt_willOverflow = (dataBusReadArea_lastCnt_willOverflowIfInc && dataBusReadArea_lastCnt_willIncrement);
  always @(*) begin
    dataBusReadArea_lastCnt_valueNext = (dataBusReadArea_lastCnt_value + _zz_dataBusReadArea_lastCnt_valueNext);
    if(dataBusReadArea_lastCnt_willClear) begin
      dataBusReadArea_lastCnt_valueNext = 32'h0;
    end
  end

  assign toplevel_pippenger_1_io_dataIn_fire = (dataBusReadArea_inputValid && pippenger_1_io_dataIn_ready);
  assign pippenger_1_io_dataIn_payload_fragment_P_X = dataBusReadArea_outputData_0[376:0];
  assign pippenger_1_io_dataIn_payload_fragment_P_Y = dataBusReadArea_outputData_1[376:0];
  assign pippenger_1_io_dataIn_payload_fragment_P_T = dataBusReadArea_outputData_2[376:0];
  assign pippenger_1_io_dataIn_payload_fragment_K = dataBusReadArea_outputData_3[252:0];
  assign dataBusReadArea_inputDMA_io_streamBus_ready = ((! dataBusReadArea_inputValid) || pippenger_1_io_dataIn_ready);
  assign toplevel_dataBusReadArea_inputDMA_io_streamBus_fire = (dataBusReadArea_inputDMA_io_streamBus_valid && dataBusReadArea_inputDMA_io_streamBus_ready);
  always @(*) begin
    dataBusWriteArea_outputCnt_willIncrement = 1'b0;
    if(io_dataBus_w_fire) begin
      dataBusWriteArea_outputCnt_willIncrement = 1'b1;
    end
  end

  assign dataBusWriteArea_outputCnt_willClear = 1'b0;
  assign dataBusWriteArea_outputCnt_willOverflow = (dataBusWriteArea_outputCnt_willOverflowIfInc && dataBusWriteArea_outputCnt_willIncrement);
  always @(*) begin
    dataBusWriteArea_outputCnt_valueNext = (dataBusWriteArea_outputCnt_value + _zz_dataBusWriteArea_outputCnt_valueNext);
    if(dataBusWriteArea_outputCnt_willClear) begin
      dataBusWriteArea_outputCnt_valueNext = 2'b00;
    end
  end

  assign dataBus_awvalid = dataBusWriteArea_addressOutputValid;
  assign dataBus_awaddr = startWriteAddress;
  assign dataBus_awlen = 8'h03;
  assign dataBus_wvalid = dataBusWriteArea_dataOutputValid;
  assign dataBus_wdata = {135'd0, _zz_dataBus_wdata};
  assign dataBus_wlast = dataBusWriteArea_outputCnt_willOverflowIfInc;
  assign io_dataBus_w_fire = (dataBus_wvalid && dataBus_wready);
  assign dataBus_bready = 1'b1;
  assign when_AxiLite4SlaveFactory_l68 = ((slaveFactory_writeAddressMasked & (~ 6'h03)) == 6'h20);
  assign when_AxiLite4SlaveFactory_l68_1 = ((slaveFactory_writeAddressMasked & (~ 6'h03)) == 6'h24);
  assign when_AxiLite4SlaveFactory_l68_2 = ((slaveFactory_writeAddressMasked & (~ 6'h03)) == 6'h28);
  assign when_AxiLite4SlaveFactory_l68_3 = ((slaveFactory_writeAddressMasked & (~ 6'h03)) == 6'h2c);
  assign when_AxiLite4SlaveFactory_l86 = ((slaveFactory_readAddressMasked & (~ 6'h03)) == 6'h20);
  assign when_AxiLite4SlaveFactory_l86_1 = ((slaveFactory_readAddressMasked & (~ 6'h03)) == 6'h24);
  assign when_AxiLite4SlaveFactory_l86_2 = ((slaveFactory_readAddressMasked & (~ 6'h03)) == 6'h28);
  assign when_AxiLite4SlaveFactory_l86_3 = ((slaveFactory_readAddressMasked & (~ 6'h03)) == 6'h2c);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      readStart <= 1'b0;
      writeStart <= 1'b0;
      _zz_s_axi_control_bvalid_1 <= 1'b0;
      io_s_axi_control_ar_rValid <= 1'b0;
      dataBusReadArea_inputCnt_value <= 2'b00;
      dataBusReadArea_inputCnt_willOverflowIfInc <= 1'b0;
      dataBusReadArea_inputValid <= 1'b0;
      dataBusReadArea_lastCnt_value <= 32'h0;
      dataBusReadArea_lastCnt_willOverflowIfInc <= 1'b0;
      dataBusWriteArea_outputCnt_value <= 2'b00;
      dataBusWriteArea_outputCnt_willOverflowIfInc <= 1'b0;
      dataBusWriteArea_dataOutputValid <= 1'b0;
      dataBusWriteArea_addressOutputValid <= 1'b0;
    end else begin
      if(startRise) begin
        readStart <= 1'b1;
      end
      if(startRise) begin
        writeStart <= 1'b1;
      end
      if(_zz_slaveFactory_writeJoinEvent_translated_ready_1) begin
        _zz_s_axi_control_bvalid_1 <= (slaveFactory_writeJoinEvent_translated_valid && _zz_slaveFactory_writeJoinEvent_translated_ready);
      end
      if(s_axi_control_arready) begin
        io_s_axi_control_ar_rValid <= s_axi_control_arvalid;
      end
      if(dataBusReadArea_inputDMA_io_done) begin
        readStart <= 1'b0;
      end
      dataBusReadArea_inputCnt_value <= dataBusReadArea_inputCnt_valueNext;
      dataBusReadArea_inputCnt_willOverflowIfInc <= (dataBusReadArea_inputCnt_valueNext == 2'b10);
      dataBusReadArea_lastCnt_value <= dataBusReadArea_lastCnt_valueNext;
      dataBusReadArea_lastCnt_willOverflowIfInc <= (dataBusReadArea_lastCnt_valueNext == 32'hffffffff);
      if(dataBusReadArea_inputCnt_willOverflow) begin
        dataBusReadArea_inputValid <= 1'b1;
      end else begin
        if(pippenger_1_io_dataIn_ready) begin
          dataBusReadArea_inputValid <= 1'b0;
        end
      end
      dataBusWriteArea_outputCnt_value <= dataBusWriteArea_outputCnt_valueNext;
      dataBusWriteArea_outputCnt_willOverflowIfInc <= (dataBusWriteArea_outputCnt_valueNext == 2'b11);
      if(pippenger_1_io_dataOut_valid) begin
        dataBusWriteArea_dataOutputValid <= 1'b1;
      end else begin
        if(dataBusWriteArea_outputCnt_willOverflow) begin
          dataBusWriteArea_dataOutputValid <= 1'b0;
        end
      end
      if(pippenger_1_io_dataOut_valid) begin
        dataBusWriteArea_addressOutputValid <= 1'b1;
      end else begin
        if(dataBus_arready) begin
          dataBusWriteArea_addressOutputValid <= 1'b0;
        end
      end
      if(dataBus_bvalid) begin
        writeStart <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    pageNum <= (_zz_pageNum + 28'h0000002);
    if(_zz_slaveFactory_writeJoinEvent_translated_ready_1) begin
      _zz_s_axi_control_bresp <= slaveFactory_writeJoinEvent_translated_payload_resp;
    end
    if(s_axi_control_arready) begin
      io_s_axi_control_ar_rData_addr <= s_axi_control_araddr;
      io_s_axi_control_ar_rData_prot <= s_axi_control_arprot;
    end
    _zz_io_dataIn_payload_last <= (dataBusReadArea_lastCnt_valueNext == {num,6'h3f});
    if(toplevel_dataBusReadArea_inputDMA_io_streamBus_fire) begin
      dataBusReadArea_inputData_0 <= dataBusReadArea_inputData_1;
      dataBusReadArea_inputData_1 <= dataBusReadArea_inputData_2;
      dataBusReadArea_inputData_2 <= dataBusReadArea_inputDMA_io_streamBus_payload;
    end
    if(pippenger_1_io_dataOut_valid) begin
      dataBusWriteArea_dataReg_0 <= pippenger_1_io_dataOut_payload_X;
      dataBusWriteArea_dataReg_1 <= pippenger_1_io_dataOut_payload_Y;
      dataBusWriteArea_dataReg_2 <= pippenger_1_io_dataOut_payload_Z;
      dataBusWriteArea_dataReg_3 <= pippenger_1_io_dataOut_payload_T;
    end else begin
      if(dataBus_wready) begin
        dataBusWriteArea_dataReg_0 <= dataBusWriteArea_dataReg_1;
        dataBusWriteArea_dataReg_1 <= dataBusWriteArea_dataReg_2;
        dataBusWriteArea_dataReg_2 <= dataBusWriteArea_dataReg_3;
      end
    end
    case(slaveFactory_writeAddressMasked)
      6'h18 : begin
        if(slaveFactory_writeOccur) begin
          num <= s_axi_control_wdata[31 : 6];
        end
      end
      default : begin
      end
    endcase
    if(when_AxiLite4SlaveFactory_l68) begin
      if(slaveFactory_writeOccur) begin
        startReadAddress[31 : 0] <= _zz_startReadAddress;
      end
    end
    if(when_AxiLite4SlaveFactory_l68_1) begin
      if(slaveFactory_writeOccur) begin
        startReadAddress[63 : 32] <= _zz_startReadAddress_2;
      end
    end
    if(when_AxiLite4SlaveFactory_l68_2) begin
      if(slaveFactory_writeOccur) begin
        startWriteAddress[31 : 0] <= _zz_startWriteAddress;
      end
    end
    if(when_AxiLite4SlaveFactory_l68_3) begin
      if(slaveFactory_writeOccur) begin
        startWriteAddress[63 : 32] <= _zz_startWriteAddress_2;
      end
    end
  end

  always @(posedge clk) begin
    _zz_1 <= (dataBusReadArea_lastCnt_valueNext == {num,6'h3f});
  end


endmodule

module Axi4PageRDMA (
  output reg          io_axi4Bus_ar_valid,
  input               io_axi4Bus_ar_ready,
  output reg [63:0]   io_axi4Bus_ar_payload_addr,
  output reg [7:0]    io_axi4Bus_ar_payload_len,
  input               io_axi4Bus_r_valid,
  output              io_axi4Bus_r_ready,
  input      [511:0]  io_axi4Bus_r_payload_data,
  input               io_axi4Bus_r_payload_last,
  output              io_streamBus_valid,
  input               io_streamBus_ready,
  output     [511:0]  io_streamBus_payload,
  input               io_work,
  input      [63:0]   io_address,
  input      [27:0]   io_pageNum,
  output reg          io_done,
  input               clk,
  input               resetn
);

  wire                readFifo_io_push_ready;
  wire                readFifo_io_pop_valid;
  wire       [511:0]  readFifo_io_pop_payload;
  wire       [7:0]    readFifo_io_pushPtr;
  wire       [7:0]    readFifo_io_popPtr;
  wire       [27:0]   _zz_readArea_addressCnt_valueNext;
  wire       [0:0]    _zz_readArea_addressCnt_valueNext_1;
  wire       [1:0]    _zz_readArea_outStandingCnt_valueNext;
  wire       [0:0]    _zz_readArea_outStandingCnt_valueNext_1;
  wire       [51:0]   _zz_io_axi4Bus_ar_payload_addr;
  wire       [51:0]   _zz_io_axi4Bus_ar_payload_addr_1;
  wire                io_axi4Bus_r_translated_valid;
  wire                io_axi4Bus_r_translated_ready;
  wire       [511:0]  io_axi4Bus_r_translated_payload;
  reg                 readArea_addressCnt_willIncrement;
  reg                 readArea_addressCnt_willClear;
  reg        [27:0]   readArea_addressCnt_valueNext;
  reg        [27:0]   readArea_addressCnt_value;
  reg                 readArea_addressCnt_willOverflowIfInc;
  wire                readArea_addressCnt_willOverflow;
  reg                 readArea_outStandingCnt_willIncrement;
  wire                readArea_outStandingCnt_willClear;
  reg        [1:0]    readArea_outStandingCnt_valueNext;
  reg        [1:0]    readArea_outStandingCnt_value;
  reg                 readArea_outStandingCnt_willOverflowIfInc;
  wire                readArea_outStandingCnt_willOverflow;
  wire       [1:0]    _zz_io_axi4Bus_ar_valid;
  reg                 _zz_io_axi4Bus_ar_valid_1;
  wire                io_axi4Bus_ar_fire;
  reg                 _zz_1;

  assign _zz_readArea_addressCnt_valueNext_1 = readArea_addressCnt_willIncrement;
  assign _zz_readArea_addressCnt_valueNext = {27'd0, _zz_readArea_addressCnt_valueNext_1};
  assign _zz_readArea_outStandingCnt_valueNext_1 = readArea_outStandingCnt_willIncrement;
  assign _zz_readArea_outStandingCnt_valueNext = {1'd0, _zz_readArea_outStandingCnt_valueNext_1};
  assign _zz_io_axi4Bus_ar_payload_addr = (io_address[63 : 12] + _zz_io_axi4Bus_ar_payload_addr_1);
  assign _zz_io_axi4Bus_ar_payload_addr_1 = {24'd0, readArea_addressCnt_value};
  FIFO readFifo (
    .io_push_valid   (io_axi4Bus_r_translated_valid         ), //i
    .io_push_ready   (readFifo_io_push_ready                ), //o
    .io_push_payload (io_axi4Bus_r_translated_payload[511:0]), //i
    .io_pop_valid    (readFifo_io_pop_valid                 ), //o
    .io_pop_ready    (io_streamBus_ready                    ), //i
    .io_pop_payload  (readFifo_io_pop_payload[511:0]        ), //o
    .io_pushPtr      (readFifo_io_pushPtr[7:0]              ), //o
    .io_popPtr       (readFifo_io_popPtr[7:0]               ), //o
    .clk             (clk                                   ), //i
    .resetn          (resetn                                )  //i
  );
  assign io_streamBus_valid = readFifo_io_pop_valid;
  assign io_streamBus_payload = readFifo_io_pop_payload;
  assign io_axi4Bus_r_translated_valid = io_axi4Bus_r_valid;
  assign io_axi4Bus_r_ready = io_axi4Bus_r_translated_ready;
  assign io_axi4Bus_r_translated_payload = io_axi4Bus_r_payload_data;
  assign io_axi4Bus_r_translated_ready = readFifo_io_push_ready;
  always @(*) begin
    readArea_addressCnt_willIncrement = 1'b0;
    if(io_axi4Bus_ar_fire) begin
      readArea_addressCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    readArea_addressCnt_willClear = 1'b0;
    if(io_axi4Bus_ar_fire) begin
      if(_zz_1) begin
        readArea_addressCnt_willClear = 1'b1;
      end
    end
  end

  assign readArea_addressCnt_willOverflow = (readArea_addressCnt_willOverflowIfInc && readArea_addressCnt_willIncrement);
  always @(*) begin
    readArea_addressCnt_valueNext = (readArea_addressCnt_value + _zz_readArea_addressCnt_valueNext);
    if(readArea_addressCnt_willClear) begin
      readArea_addressCnt_valueNext = 28'h0;
    end
  end

  always @(*) begin
    readArea_outStandingCnt_willIncrement = 1'b0;
    if(io_axi4Bus_ar_fire) begin
      readArea_outStandingCnt_willIncrement = 1'b1;
    end
  end

  assign readArea_outStandingCnt_willClear = 1'b0;
  assign readArea_outStandingCnt_willOverflow = (readArea_outStandingCnt_willOverflowIfInc && readArea_outStandingCnt_willIncrement);
  always @(*) begin
    readArea_outStandingCnt_valueNext = (readArea_outStandingCnt_value + _zz_readArea_outStandingCnt_valueNext);
    if(readArea_outStandingCnt_willClear) begin
      readArea_outStandingCnt_valueNext = 2'b00;
    end
  end

  always @(*) begin
    io_axi4Bus_ar_valid = 1'b0;
    if(io_work) begin
      io_axi4Bus_ar_valid = _zz_io_axi4Bus_ar_valid_1;
    end
  end

  always @(*) begin
    io_axi4Bus_ar_payload_addr = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(io_work) begin
      io_axi4Bus_ar_payload_addr = {_zz_io_axi4Bus_ar_payload_addr,12'h0};
    end
  end

  always @(*) begin
    io_axi4Bus_ar_payload_len = 8'bxxxxxxxx;
    if(io_work) begin
      io_axi4Bus_ar_payload_len = 8'h3f;
    end
  end

  always @(*) begin
    io_done = 1'b0;
    if(io_axi4Bus_ar_fire) begin
      if(_zz_1) begin
        io_done = 1'b1;
      end
    end
  end

  assign _zz_io_axi4Bus_ar_valid = readFifo_io_popPtr[7 : 6];
  assign io_axi4Bus_ar_fire = (io_axi4Bus_ar_valid && io_axi4Bus_ar_ready);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      readArea_addressCnt_value <= 28'h0;
      readArea_addressCnt_willOverflowIfInc <= 1'b0;
      readArea_outStandingCnt_value <= 2'b00;
      readArea_outStandingCnt_willOverflowIfInc <= 1'b0;
    end else begin
      readArea_addressCnt_value <= readArea_addressCnt_valueNext;
      readArea_addressCnt_willOverflowIfInc <= (readArea_addressCnt_valueNext == 28'hfffffff);
      readArea_outStandingCnt_value <= readArea_outStandingCnt_valueNext;
      readArea_outStandingCnt_willOverflowIfInc <= (readArea_outStandingCnt_valueNext == 2'b11);
    end
  end

  always @(posedge clk) begin
    _zz_io_axi4Bus_ar_valid_1 <= (! ((readArea_outStandingCnt_valueNext[1] != _zz_io_axi4Bus_ar_valid[1]) && (readArea_outStandingCnt_valueNext[0 : 0] == _zz_io_axi4Bus_ar_valid[0 : 0])));
  end

  always @(posedge clk) begin
    _zz_1 <= (readArea_addressCnt_valueNext == io_pageNum);
  end


endmodule

module PippengerWithPAdd (
  input               io_dataIn_valid,
  output              io_dataIn_ready,
  input               io_dataIn_payload_last,
  input      [376:0]  io_dataIn_payload_fragment_P_X,
  input      [376:0]  io_dataIn_payload_fragment_P_Y,
  input      [376:0]  io_dataIn_payload_fragment_P_Z,
  input      [376:0]  io_dataIn_payload_fragment_P_T,
  input      [252:0]  io_dataIn_payload_fragment_K,
  output              io_dataOut_valid,
  input               io_dataOut_ready,
  output     [376:0]  io_dataOut_payload_X,
  output     [376:0]  io_dataOut_payload_Y,
  output     [376:0]  io_dataOut_payload_Z,
  output     [376:0]  io_dataOut_payload_T,
  input               clk,
  input               resetn
);

  wire       [376:0]  adder_0_io_s_X;
  wire       [376:0]  adder_0_io_s_Y;
  wire       [376:0]  adder_0_io_s_Z;
  wire       [376:0]  adder_0_io_s_T;
  wire       [376:0]  neg_io_n_X;
  wire       [376:0]  neg_io_n_Y;
  wire       [376:0]  neg_io_n_Z;
  wire       [376:0]  neg_io_n_T;
  wire                pippenger_1_io_dataIn_ready;
  wire                pippenger_1_io_dataOut_valid;
  wire       [376:0]  pippenger_1_io_dataOut_payload_X;
  wire       [376:0]  pippenger_1_io_dataOut_payload_Y;
  wire       [376:0]  pippenger_1_io_dataOut_payload_Z;
  wire       [376:0]  pippenger_1_io_dataOut_payload_T;
  wire       [376:0]  pippenger_1_pAddPort_0_a_X;
  wire       [376:0]  pippenger_1_pAddPort_0_a_Y;
  wire       [376:0]  pippenger_1_pAddPort_0_a_Z;
  wire       [376:0]  pippenger_1_pAddPort_0_a_T;
  wire       [376:0]  pippenger_1_pAddPort_0_b_X;
  wire       [376:0]  pippenger_1_pAddPort_0_b_Y;
  wire       [376:0]  pippenger_1_pAddPort_0_b_Z;
  wire       [376:0]  pippenger_1_pAddPort_0_b_T;
  wire       [376:0]  pippenger_1_pNegPort_a_X;
  wire       [376:0]  pippenger_1_pNegPort_a_Y;
  wire       [376:0]  pippenger_1_pNegPort_a_Z;
  wire       [376:0]  pippenger_1_pNegPort_a_T;

  PAdd adder_0 (
    .io_a_X (pippenger_1_pAddPort_0_a_X[376:0]), //i
    .io_a_Y (pippenger_1_pAddPort_0_a_Y[376:0]), //i
    .io_a_Z (pippenger_1_pAddPort_0_a_Z[376:0]), //i
    .io_a_T (pippenger_1_pAddPort_0_a_T[376:0]), //i
    .io_b_X (pippenger_1_pAddPort_0_b_X[376:0]), //i
    .io_b_Y (pippenger_1_pAddPort_0_b_Y[376:0]), //i
    .io_b_Z (pippenger_1_pAddPort_0_b_Z[376:0]), //i
    .io_b_T (pippenger_1_pAddPort_0_b_T[376:0]), //i
    .io_s_X (adder_0_io_s_X[376:0]            ), //o
    .io_s_Y (adder_0_io_s_Y[376:0]            ), //o
    .io_s_Z (adder_0_io_s_Z[376:0]            ), //o
    .io_s_T (adder_0_io_s_T[376:0]            ), //o
    .clk    (clk                              ), //i
    .resetn (resetn                           )  //i
  );
  PNeg neg (
    .io_a_X (pippenger_1_pNegPort_a_X[376:0]), //i
    .io_a_Y (pippenger_1_pNegPort_a_Y[376:0]), //i
    .io_a_Z (pippenger_1_pNegPort_a_Z[376:0]), //i
    .io_a_T (pippenger_1_pNegPort_a_T[376:0]), //i
    .io_n_X (neg_io_n_X[376:0]              ), //o
    .io_n_Y (neg_io_n_Y[376:0]              ), //o
    .io_n_Z (neg_io_n_Z[376:0]              ), //o
    .io_n_T (neg_io_n_T[376:0]              ), //o
    .clk    (clk                            ), //i
    .resetn (resetn                         )  //i
  );
  Pippenger pippenger_1 (
    .io_dataIn_valid                (io_dataIn_valid                                                                                     ), //i
    .io_dataIn_ready                (pippenger_1_io_dataIn_ready                                                                         ), //o
    .io_dataIn_payload_last         (io_dataIn_payload_last                                                                              ), //i
    .io_dataIn_payload_fragment_P_X (io_dataIn_payload_fragment_P_X[376:0]                                                               ), //i
    .io_dataIn_payload_fragment_P_Y (io_dataIn_payload_fragment_P_Y[376:0]                                                               ), //i
    .io_dataIn_payload_fragment_P_Z (io_dataIn_payload_fragment_P_Z[376:0]                                                               ), //i
    .io_dataIn_payload_fragment_P_T (io_dataIn_payload_fragment_P_T[376:0]                                                               ), //i
    .io_dataIn_payload_fragment_K   (io_dataIn_payload_fragment_K[252:0]                                                                 ), //i
    .io_dataOut_valid               (pippenger_1_io_dataOut_valid                                                                        ), //o
    .io_dataOut_ready               (io_dataOut_ready                                                                                    ), //i
    .io_dataOut_payload_X           (pippenger_1_io_dataOut_payload_X[376:0]                                                             ), //o
    .io_dataOut_payload_Y           (pippenger_1_io_dataOut_payload_Y[376:0]                                                             ), //o
    .io_dataOut_payload_Z           (pippenger_1_io_dataOut_payload_Z[376:0]                                                             ), //o
    .io_dataOut_payload_T           (pippenger_1_io_dataOut_payload_T[376:0]                                                             ), //o
    .io_pInit_X                     (377'h0                                                                                              ), //i
    .io_pInit_Y                     (377'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001), //i
    .io_pInit_Z                     (377'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001), //i
    .io_pInit_T                     (377'h0                                                                                              ), //i
    .pAddPort_0_a_X                 (pippenger_1_pAddPort_0_a_X[376:0]                                                                   ), //o
    .pAddPort_0_a_Y                 (pippenger_1_pAddPort_0_a_Y[376:0]                                                                   ), //o
    .pAddPort_0_a_Z                 (pippenger_1_pAddPort_0_a_Z[376:0]                                                                   ), //o
    .pAddPort_0_a_T                 (pippenger_1_pAddPort_0_a_T[376:0]                                                                   ), //o
    .pAddPort_0_b_X                 (pippenger_1_pAddPort_0_b_X[376:0]                                                                   ), //o
    .pAddPort_0_b_Y                 (pippenger_1_pAddPort_0_b_Y[376:0]                                                                   ), //o
    .pAddPort_0_b_Z                 (pippenger_1_pAddPort_0_b_Z[376:0]                                                                   ), //o
    .pAddPort_0_b_T                 (pippenger_1_pAddPort_0_b_T[376:0]                                                                   ), //o
    .pAddPort_0_s_X                 (adder_0_io_s_X[376:0]                                                                               ), //i
    .pAddPort_0_s_Y                 (adder_0_io_s_Y[376:0]                                                                               ), //i
    .pAddPort_0_s_Z                 (adder_0_io_s_Z[376:0]                                                                               ), //i
    .pAddPort_0_s_T                 (adder_0_io_s_T[376:0]                                                                               ), //i
    .pNegPort_a_X                   (pippenger_1_pNegPort_a_X[376:0]                                                                     ), //o
    .pNegPort_a_Y                   (pippenger_1_pNegPort_a_Y[376:0]                                                                     ), //o
    .pNegPort_a_Z                   (pippenger_1_pNegPort_a_Z[376:0]                                                                     ), //o
    .pNegPort_a_T                   (pippenger_1_pNegPort_a_T[376:0]                                                                     ), //o
    .pNegPort_n_X                   (neg_io_n_X[376:0]                                                                                   ), //i
    .pNegPort_n_Y                   (neg_io_n_Y[376:0]                                                                                   ), //i
    .pNegPort_n_Z                   (neg_io_n_Z[376:0]                                                                                   ), //i
    .pNegPort_n_T                   (neg_io_n_T[376:0]                                                                                   ), //i
    .clk                            (clk                                                                                                 ), //i
    .resetn                         (resetn                                                                                              )  //i
  );
  assign io_dataIn_ready = pippenger_1_io_dataIn_ready;
  assign io_dataOut_valid = pippenger_1_io_dataOut_valid;
  assign io_dataOut_payload_X = pippenger_1_io_dataOut_payload_X;
  assign io_dataOut_payload_Y = pippenger_1_io_dataOut_payload_Y;
  assign io_dataOut_payload_Z = pippenger_1_io_dataOut_payload_Z;
  assign io_dataOut_payload_T = pippenger_1_io_dataOut_payload_T;

endmodule

module FIFO (
  input               io_push_valid,
  output              io_push_ready,
  input      [511:0]  io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [511:0]  io_pop_payload,
  output     [7:0]    io_pushPtr,
  output     [7:0]    io_popPtr,
  input               clk,
  input               resetn
);

  reg        [511:0]  _zz_useRam_ram_port1;
  wire       [7:0]    _zz_useRam_pushPtr_valueNext;
  wire       [0:0]    _zz_useRam_pushPtr_valueNext_1;
  wire       [7:0]    _zz_useRam_popPtr_valueNext;
  wire       [0:0]    _zz_useRam_popPtr_valueNext_1;
  wire       [6:0]    _zz_useRam_ram_port;
  wire       [6:0]    _zz_useRam_ram_port_1;
  wire                _zz_useRam_ram_port_2;
  wire       [6:0]    _zz_io_pop_payload_1;
  wire                _zz_io_pop_payload_2;
  reg                 _zz_1;
  reg                 useRam_pushPtr_willIncrement;
  wire                useRam_pushPtr_willClear;
  reg        [7:0]    useRam_pushPtr_valueNext;
  reg        [7:0]    useRam_pushPtr_value;
  reg                 useRam_pushPtr_willOverflowIfInc;
  wire                useRam_pushPtr_willOverflow;
  reg                 useRam_popPtr_willIncrement;
  wire                useRam_popPtr_willClear;
  reg        [7:0]    useRam_popPtr_valueNext;
  reg        [7:0]    useRam_popPtr_value;
  reg                 useRam_popPtr_willOverflowIfInc;
  wire                useRam_popPtr_willOverflow;
  reg                 _zz_io_push_ready;
  wire                io_push_fire;
  reg                 _zz_io_pop_valid;
  wire       [7:0]    _zz_io_pop_payload;
  wire                io_pop_fire;
  reg [511:0] useRam_ram [0:127];

  assign _zz_useRam_pushPtr_valueNext_1 = useRam_pushPtr_willIncrement;
  assign _zz_useRam_pushPtr_valueNext = {7'd0, _zz_useRam_pushPtr_valueNext_1};
  assign _zz_useRam_popPtr_valueNext_1 = useRam_popPtr_willIncrement;
  assign _zz_useRam_popPtr_valueNext = {7'd0, _zz_useRam_popPtr_valueNext_1};
  assign _zz_useRam_ram_port = useRam_pushPtr_value[6:0];
  assign _zz_io_pop_payload_1 = _zz_io_pop_payload[6:0];
  assign _zz_io_pop_payload_2 = 1'b1;
  always @(posedge clk) begin
    if(_zz_1) begin
      useRam_ram[_zz_useRam_ram_port] <= io_push_payload;
    end
  end

  always @(posedge clk) begin
    if(_zz_io_pop_payload_2) begin
      _zz_useRam_ram_port1 <= useRam_ram[_zz_io_pop_payload_1];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    useRam_pushPtr_willIncrement = 1'b0;
    if(io_push_fire) begin
      useRam_pushPtr_willIncrement = 1'b1;
    end
  end

  assign useRam_pushPtr_willClear = 1'b0;
  assign useRam_pushPtr_willOverflow = (useRam_pushPtr_willOverflowIfInc && useRam_pushPtr_willIncrement);
  always @(*) begin
    useRam_pushPtr_valueNext = (useRam_pushPtr_value + _zz_useRam_pushPtr_valueNext);
    if(useRam_pushPtr_willClear) begin
      useRam_pushPtr_valueNext = 8'h0;
    end
  end

  always @(*) begin
    useRam_popPtr_willIncrement = 1'b0;
    if(io_pop_fire) begin
      useRam_popPtr_willIncrement = 1'b1;
    end
  end

  assign useRam_popPtr_willClear = 1'b0;
  assign useRam_popPtr_willOverflow = (useRam_popPtr_willOverflowIfInc && useRam_popPtr_willIncrement);
  always @(*) begin
    useRam_popPtr_valueNext = (useRam_popPtr_value + _zz_useRam_popPtr_valueNext);
    if(useRam_popPtr_willClear) begin
      useRam_popPtr_valueNext = 8'h0;
    end
  end

  assign io_pushPtr = useRam_pushPtr_value;
  assign io_popPtr = useRam_popPtr_value;
  assign io_push_ready = _zz_io_push_ready;
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign io_pop_valid = _zz_io_pop_valid;
  assign _zz_io_pop_payload = useRam_popPtr_valueNext;
  assign io_pop_payload = _zz_useRam_ram_port1;
  assign io_pop_fire = (io_pop_valid && io_pop_ready);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      useRam_pushPtr_value <= 8'h0;
      useRam_pushPtr_willOverflowIfInc <= 1'b0;
      useRam_popPtr_value <= 8'h0;
      useRam_popPtr_willOverflowIfInc <= 1'b0;
      _zz_io_push_ready <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      useRam_pushPtr_value <= useRam_pushPtr_valueNext;
      useRam_pushPtr_willOverflowIfInc <= (useRam_pushPtr_valueNext == 8'hff);
      useRam_popPtr_value <= useRam_popPtr_valueNext;
      useRam_popPtr_willOverflowIfInc <= (useRam_popPtr_valueNext == 8'hff);
      _zz_io_push_ready <= (! ((useRam_pushPtr_valueNext[7] != useRam_popPtr_value[7]) && (useRam_pushPtr_valueNext[6 : 0] == useRam_popPtr_value[6 : 0])));
      _zz_io_pop_valid <= (! (useRam_pushPtr_value == useRam_popPtr_valueNext));
    end
  end


endmodule

module Pippenger (
  input               io_dataIn_valid,
  output              io_dataIn_ready,
  input               io_dataIn_payload_last,
  input      [376:0]  io_dataIn_payload_fragment_P_X,
  input      [376:0]  io_dataIn_payload_fragment_P_Y,
  input      [376:0]  io_dataIn_payload_fragment_P_Z,
  input      [376:0]  io_dataIn_payload_fragment_P_T,
  input      [252:0]  io_dataIn_payload_fragment_K,
  output              io_dataOut_valid,
  input               io_dataOut_ready,
  output     [376:0]  io_dataOut_payload_X,
  output     [376:0]  io_dataOut_payload_Y,
  output     [376:0]  io_dataOut_payload_Z,
  output     [376:0]  io_dataOut_payload_T,
  input      [376:0]  io_pInit_X,
  input      [376:0]  io_pInit_Y,
  input      [376:0]  io_pInit_Z,
  input      [376:0]  io_pInit_T,
  output     [376:0]  pAddPort_0_a_X,
  output     [376:0]  pAddPort_0_a_Y,
  output     [376:0]  pAddPort_0_a_Z,
  output     [376:0]  pAddPort_0_a_T,
  output     [376:0]  pAddPort_0_b_X,
  output     [376:0]  pAddPort_0_b_Y,
  output     [376:0]  pAddPort_0_b_Z,
  output     [376:0]  pAddPort_0_b_T,
  input      [376:0]  pAddPort_0_s_X,
  input      [376:0]  pAddPort_0_s_Y,
  input      [376:0]  pAddPort_0_s_Z,
  input      [376:0]  pAddPort_0_s_T,
  output     [376:0]  pNegPort_a_X,
  output     [376:0]  pNegPort_a_Y,
  output     [376:0]  pNegPort_a_Z,
  output     [376:0]  pNegPort_a_T,
  input      [376:0]  pNegPort_n_X,
  input      [376:0]  pNegPort_n_Y,
  input      [376:0]  pNegPort_n_Z,
  input      [376:0]  pNegPort_n_T,
  input               clk,
  input               resetn
);
  localparam fsm_enumDef_flushing = 4'd1;
  localparam fsm_enumDef_stage1 = 4'd2;
  localparam fsm_enumDef_stage2 = 4'd4;
  localparam fsm_enumDef_stage3 = 4'd8;

  reg                 stateRam_0_io_we_0;
  reg                 stateRam_0_io_we_1;
  reg        [16:0]   stateRam_0_io_address_0;
  reg        [16:0]   stateRam_0_io_address_1;
  reg                 stateRam_0_io_flush;
  reg        [16:0]   stateRam_0_io_flushCnt;
  reg                 dataRam_0_io_we_0;
  reg                 dataRam_0_io_we_1;
  reg        [16:0]   dataRam_0_io_address_0;
  reg        [16:0]   dataRam_0_io_address_1;
  reg        [376:0]  dataRam_0_io_wData_0_X;
  reg        [376:0]  dataRam_0_io_wData_0_Y;
  reg        [376:0]  dataRam_0_io_wData_0_Z;
  reg        [376:0]  dataRam_0_io_wData_0_T;
  reg        [376:0]  dataRam_0_io_wData_1_X;
  reg        [376:0]  dataRam_0_io_wData_1_Y;
  reg        [376:0]  dataRam_0_io_wData_1_Z;
  reg        [376:0]  dataRam_0_io_wData_1_T;
  reg                 dataRam_0_io_state_1;
  reg                 fifo_0_io_dataIn_0_valid;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_a_X;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_a_Y;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_a_Z;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_a_T;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_b_X;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_b_Y;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_b_Z;
  reg        [376:0]  fifo_0_io_dataIn_0_payload_b_T;
  reg        [16:0]   fifo_0_io_dataIn_0_payload_address;
  reg                 fifo_0_io_dataIn_1_valid;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_a_X;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_a_Y;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_a_Z;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_a_T;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_b_X;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_b_Y;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_b_Z;
  reg        [376:0]  fifo_0_io_dataIn_1_payload_b_T;
  reg        [16:0]   fifo_0_io_dataIn_1_payload_address;
  wire                stateRam_0_io_state_0;
  wire                stateRam_0_io_state_1;
  wire       [376:0]  dataRam_0_io_rData_0_X;
  wire       [376:0]  dataRam_0_io_rData_0_Y;
  wire       [376:0]  dataRam_0_io_rData_0_Z;
  wire       [376:0]  dataRam_0_io_rData_0_T;
  wire       [376:0]  dataRam_0_io_rData_1_X;
  wire       [376:0]  dataRam_0_io_rData_1_Y;
  wire       [376:0]  dataRam_0_io_rData_1_Z;
  wire       [376:0]  dataRam_0_io_rData_1_T;
  wire                fifo_0_io_dataOut_valid;
  wire       [376:0]  fifo_0_io_dataOut_payload_a_X;
  wire       [376:0]  fifo_0_io_dataOut_payload_a_Y;
  wire       [376:0]  fifo_0_io_dataOut_payload_a_Z;
  wire       [376:0]  fifo_0_io_dataOut_payload_a_T;
  wire       [376:0]  fifo_0_io_dataOut_payload_b_X;
  wire       [376:0]  fifo_0_io_dataOut_payload_b_Y;
  wire       [376:0]  fifo_0_io_dataOut_payload_b_Z;
  wire       [376:0]  fifo_0_io_dataOut_payload_b_T;
  wire       [16:0]   fifo_0_io_dataOut_payload_address;
  wire       [239:0]  _zz_dataInBuffer_dataReg_fragment_K;
  wire       [16:0]   _zz_flushing_flushCnt_valueNext;
  wire       [0:0]    _zz_flushing_flushCnt_valueNext_1;
  wire       [31:0]   _zz_stage1_NCnt_valueNext;
  wire       [0:0]    _zz_stage1_NCnt_valueNext_1;
  wire       [4:0]    _zz_stage1_GCnt_valueNext;
  wire       [0:0]    _zz_stage1_GCnt_valueNext_1;
  wire       [8:0]    _zz_stage1_emptyCnt_valueNext;
  wire       [0:0]    _zz_stage1_emptyCnt_valueNext_1;
  wire       [12:0]   _zz_stage1_inputBarrelID_0;
  wire       [13:0]   _zz_stage1_inputBarrelID_0_1;
  wire       [1:0]    _zz_stage1_inputBarrelID_0_2;
  wire       [12:0]   _zz__zz_stage1_inputBarrelIDAbs_0;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0_1;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0_2;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0_3;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0_4;
  wire       [0:0]    _zz_stage1_inputBarrelIDAbs_0_5;
  wire       [12:0]   _zz__zz_stage1_inputValid_0;
  wire       [11:0]   _zz_stage2_wCnt_valueNext;
  wire       [0:0]    _zz_stage2_wCnt_valueNext_1;
  wire       [4:0]    _zz_stage2_GCnt_valueNext;
  wire       [0:0]    _zz_stage2_GCnt_valueNext_1;
  wire       [1:0]    _zz_stage2_calCnt_valueNext;
  wire       [0:0]    _zz_stage2_calCnt_valueNext_1;
  wire       [8:0]    _zz_stage2_waitCnt_valueNext;
  wire       [0:0]    _zz_stage2_waitCnt_valueNext_1;
  wire       [4:0]    _zz_stage3_GCnt_valueNext;
  wire       [0:0]    _zz_stage3_GCnt_valueNext_1;
  wire       [3:0]    _zz_stage3_doubleCnt_valueNext;
  wire       [0:0]    _zz_stage3_doubleCnt_valueNext_1;
  wire       [8:0]    _zz_stage3_doubleWaitCnt_valueNext;
  wire       [0:0]    _zz_stage3_doubleWaitCnt_valueNext_1;
  wire       [8:0]    _zz_stage3_addWaitCnt_valueNext;
  wire       [0:0]    _zz_stage3_addWaitCnt_valueNext_1;
  wire       [11:0]   _zz_io_address_0;
  wire       [11:0]   _zz_io_address_0_1;
  wire       [11:0]   _zz_io_address_0_2;
  wire       [11:0]   _zz_io_address_1;
  wire       [11:0]   _zz_io_address_1_1;
  wire       [11:0]   _zz_io_address_1_2;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address_1;
  wire       [11:0]   _zz__zz_io_dataIn_1_payload_address_2;
  wire       [4:0]    _zz_io_address_1_3;
  wire       [4:0]    _zz_io_address_1_4;
  wire       [0:0]    _zz_io_address_1_5;
  wire       [4:0]    _zz__zz_io_dataIn_1_payload_address_30;
  wire       [0:0]    _zz__zz_io_dataIn_1_payload_address_30_1;
  wire                dataInBuffer_bufferOut_valid;
  reg                 dataInBuffer_bufferOut_ready;
  wire                dataInBuffer_bufferOut_payload_last;
  wire       [376:0]  dataInBuffer_bufferOut_payload_fragment_P_X;
  wire       [376:0]  dataInBuffer_bufferOut_payload_fragment_P_Y;
  wire       [376:0]  dataInBuffer_bufferOut_payload_fragment_P_Z;
  wire       [376:0]  dataInBuffer_bufferOut_payload_fragment_P_T;
  wire       [252:0]  dataInBuffer_bufferOut_payload_fragment_K;
  reg                 dataInBuffer_shift;
  reg                 dataInBuffer_validReg;
  reg                 dataInBuffer_dataReg_last;
  reg        [376:0]  dataInBuffer_dataReg_fragment_P_X;
  reg        [376:0]  dataInBuffer_dataReg_fragment_P_Y;
  reg        [376:0]  dataInBuffer_dataReg_fragment_P_Z;
  reg        [376:0]  dataInBuffer_dataReg_fragment_P_T;
  reg        [252:0]  dataInBuffer_dataReg_fragment_K;
  wire                shiftRegs_validIn_0;
  wire       [16:0]   shiftRegs_addressIn_0;
  reg                 shiftRegs_validIn_delay_1_0;
  reg                 shiftRegs_validIn_delay_2_0;
  reg                 shiftRegs_validIn_delay_3_0;
  reg                 shiftRegs_validIn_delay_4_0;
  reg                 shiftRegs_validIn_delay_5_0;
  reg                 shiftRegs_validIn_delay_6_0;
  reg                 shiftRegs_validIn_delay_7_0;
  reg                 shiftRegs_validIn_delay_8_0;
  reg                 shiftRegs_validIn_delay_9_0;
  reg                 shiftRegs_validIn_delay_10_0;
  reg                 shiftRegs_validIn_delay_11_0;
  reg                 shiftRegs_validIn_delay_12_0;
  reg                 shiftRegs_validIn_delay_13_0;
  reg                 shiftRegs_validIn_delay_14_0;
  reg                 shiftRegs_validIn_delay_15_0;
  reg                 shiftRegs_validIn_delay_16_0;
  reg                 shiftRegs_validIn_delay_17_0;
  reg                 shiftRegs_validIn_delay_18_0;
  reg                 shiftRegs_validIn_delay_19_0;
  reg                 shiftRegs_validIn_delay_20_0;
  reg                 shiftRegs_validIn_delay_21_0;
  reg                 shiftRegs_validIn_delay_22_0;
  reg                 shiftRegs_validIn_delay_23_0;
  reg                 shiftRegs_validIn_delay_24_0;
  reg                 shiftRegs_validIn_delay_25_0;
  reg                 shiftRegs_validIn_delay_26_0;
  reg                 shiftRegs_validIn_delay_27_0;
  reg                 shiftRegs_validIn_delay_28_0;
  reg                 shiftRegs_validIn_delay_29_0;
  reg                 shiftRegs_validIn_delay_30_0;
  reg                 shiftRegs_validIn_delay_31_0;
  reg                 shiftRegs_validIn_delay_32_0;
  reg                 shiftRegs_validIn_delay_33_0;
  reg                 shiftRegs_validIn_delay_34_0;
  reg                 shiftRegs_validIn_delay_35_0;
  reg                 shiftRegs_validIn_delay_36_0;
  reg                 shiftRegs_validIn_delay_37_0;
  reg                 shiftRegs_validIn_delay_38_0;
  reg                 shiftRegs_validIn_delay_39_0;
  reg                 shiftRegs_validIn_delay_40_0;
  reg                 shiftRegs_validIn_delay_41_0;
  reg                 shiftRegs_validIn_delay_42_0;
  reg                 shiftRegs_validIn_delay_43_0;
  reg                 shiftRegs_validIn_delay_44_0;
  reg                 shiftRegs_validIn_delay_45_0;
  reg                 shiftRegs_validIn_delay_46_0;
  reg                 shiftRegs_validIn_delay_47_0;
  reg                 shiftRegs_validIn_delay_48_0;
  reg                 shiftRegs_validIn_delay_49_0;
  reg                 shiftRegs_validIn_delay_50_0;
  reg                 shiftRegs_validIn_delay_51_0;
  reg                 shiftRegs_validIn_delay_52_0;
  reg                 shiftRegs_validIn_delay_53_0;
  reg                 shiftRegs_validIn_delay_54_0;
  reg                 shiftRegs_validIn_delay_55_0;
  reg                 shiftRegs_validIn_delay_56_0;
  reg                 shiftRegs_validIn_delay_57_0;
  reg                 shiftRegs_validIn_delay_58_0;
  reg                 shiftRegs_validIn_delay_59_0;
  reg                 shiftRegs_validIn_delay_60_0;
  reg                 shiftRegs_validIn_delay_61_0;
  reg                 shiftRegs_validIn_delay_62_0;
  reg                 shiftRegs_validIn_delay_63_0;
  reg                 shiftRegs_validIn_delay_64_0;
  reg                 shiftRegs_validIn_delay_65_0;
  reg                 shiftRegs_validIn_delay_66_0;
  reg                 shiftRegs_validIn_delay_67_0;
  reg                 shiftRegs_validIn_delay_68_0;
  reg                 shiftRegs_validIn_delay_69_0;
  reg                 shiftRegs_validIn_delay_70_0;
  reg                 shiftRegs_validIn_delay_71_0;
  reg                 shiftRegs_validIn_delay_72_0;
  reg                 shiftRegs_validIn_delay_73_0;
  reg                 shiftRegs_validIn_delay_74_0;
  reg                 shiftRegs_validIn_delay_75_0;
  reg                 shiftRegs_validIn_delay_76_0;
  reg                 shiftRegs_validIn_delay_77_0;
  reg                 shiftRegs_validIn_delay_78_0;
  reg                 shiftRegs_validIn_delay_79_0;
  reg                 shiftRegs_validIn_delay_80_0;
  reg                 shiftRegs_validIn_delay_81_0;
  reg                 shiftRegs_validIn_delay_82_0;
  reg                 shiftRegs_validIn_delay_83_0;
  reg                 shiftRegs_validIn_delay_84_0;
  reg                 shiftRegs_validIn_delay_85_0;
  reg                 shiftRegs_validIn_delay_86_0;
  reg                 shiftRegs_validIn_delay_87_0;
  reg                 shiftRegs_validIn_delay_88_0;
  reg                 shiftRegs_validIn_delay_89_0;
  reg                 shiftRegs_validIn_delay_90_0;
  reg                 shiftRegs_validIn_delay_91_0;
  reg                 shiftRegs_validIn_delay_92_0;
  reg                 shiftRegs_validIn_delay_93_0;
  reg                 shiftRegs_validIn_delay_94_0;
  reg                 shiftRegs_validIn_delay_95_0;
  reg                 shiftRegs_validIn_delay_96_0;
  reg                 shiftRegs_validIn_delay_97_0;
  reg                 shiftRegs_validIn_delay_98_0;
  reg                 shiftRegs_validIn_delay_99_0;
  reg                 shiftRegs_validIn_delay_100_0;
  reg                 shiftRegs_validIn_delay_101_0;
  reg                 shiftRegs_validIn_delay_102_0;
  reg                 shiftRegs_validIn_delay_103_0;
  reg                 shiftRegs_validIn_delay_104_0;
  reg                 shiftRegs_validIn_delay_105_0;
  reg                 shiftRegs_validIn_delay_106_0;
  reg                 shiftRegs_validIn_delay_107_0;
  reg                 shiftRegs_validIn_delay_108_0;
  reg                 shiftRegs_validIn_delay_109_0;
  reg                 shiftRegs_validIn_delay_110_0;
  reg                 shiftRegs_validIn_delay_111_0;
  reg                 shiftRegs_validIn_delay_112_0;
  reg                 shiftRegs_validIn_delay_113_0;
  reg                 shiftRegs_validIn_delay_114_0;
  reg                 shiftRegs_validIn_delay_115_0;
  reg                 shiftRegs_validIn_delay_116_0;
  reg                 shiftRegs_validIn_delay_117_0;
  reg                 shiftRegs_validIn_delay_118_0;
  reg                 shiftRegs_validIn_delay_119_0;
  reg                 shiftRegs_validIn_delay_120_0;
  reg                 shiftRegs_validIn_delay_121_0;
  reg                 shiftRegs_validIn_delay_122_0;
  reg                 shiftRegs_validIn_delay_123_0;
  reg                 shiftRegs_validIn_delay_124_0;
  reg                 shiftRegs_validIn_delay_125_0;
  reg                 shiftRegs_validIn_delay_126_0;
  reg                 shiftRegs_validIn_delay_127_0;
  reg                 shiftRegs_validIn_delay_128_0;
  reg                 shiftRegs_validIn_delay_129_0;
  reg                 shiftRegs_validIn_delay_130_0;
  reg                 shiftRegs_validIn_delay_131_0;
  reg                 shiftRegs_validIn_delay_132_0;
  reg                 shiftRegs_validIn_delay_133_0;
  reg                 shiftRegs_validIn_delay_134_0;
  reg                 shiftRegs_validIn_delay_135_0;
  reg                 shiftRegs_validIn_delay_136_0;
  reg                 shiftRegs_validIn_delay_137_0;
  reg                 shiftRegs_validIn_delay_138_0;
  reg                 shiftRegs_validIn_delay_139_0;
  reg                 shiftRegs_validIn_delay_140_0;
  reg                 shiftRegs_validIn_delay_141_0;
  reg                 shiftRegs_validIn_delay_142_0;
  reg                 shiftRegs_validIn_delay_143_0;
  reg                 shiftRegs_validIn_delay_144_0;
  reg                 shiftRegs_validIn_delay_145_0;
  reg                 shiftRegs_validIn_delay_146_0;
  reg                 shiftRegs_validIn_delay_147_0;
  reg                 shiftRegs_validIn_delay_148_0;
  reg                 shiftRegs_validIn_delay_149_0;
  reg                 shiftRegs_validIn_delay_150_0;
  reg                 shiftRegs_validIn_delay_151_0;
  reg                 shiftRegs_validIn_delay_152_0;
  reg                 shiftRegs_validIn_delay_153_0;
  reg                 shiftRegs_validIn_delay_154_0;
  reg                 shiftRegs_validIn_delay_155_0;
  reg                 shiftRegs_validIn_delay_156_0;
  reg                 shiftRegs_validIn_delay_157_0;
  reg                 shiftRegs_validIn_delay_158_0;
  reg                 shiftRegs_validIn_delay_159_0;
  reg                 shiftRegs_validIn_delay_160_0;
  reg                 shiftRegs_validIn_delay_161_0;
  reg                 shiftRegs_validIn_delay_162_0;
  reg                 shiftRegs_validIn_delay_163_0;
  reg                 shiftRegs_validIn_delay_164_0;
  reg                 shiftRegs_validIn_delay_165_0;
  reg                 shiftRegs_validIn_delay_166_0;
  reg                 shiftRegs_validIn_delay_167_0;
  reg                 shiftRegs_validIn_delay_168_0;
  reg                 shiftRegs_validIn_delay_169_0;
  reg                 shiftRegs_validIn_delay_170_0;
  reg                 shiftRegs_validIn_delay_171_0;
  reg                 shiftRegs_validIn_delay_172_0;
  reg                 shiftRegs_validIn_delay_173_0;
  reg                 shiftRegs_validIn_delay_174_0;
  reg                 shiftRegs_validIn_delay_175_0;
  reg                 shiftRegs_validIn_delay_176_0;
  reg                 shiftRegs_validIn_delay_177_0;
  reg                 shiftRegs_validIn_delay_178_0;
  reg                 shiftRegs_validIn_delay_179_0;
  reg                 shiftRegs_validIn_delay_180_0;
  reg                 shiftRegs_validIn_delay_181_0;
  reg                 shiftRegs_validIn_delay_182_0;
  reg                 shiftRegs_validIn_delay_183_0;
  reg                 shiftRegs_validIn_delay_184_0;
  reg                 shiftRegs_validIn_delay_185_0;
  reg                 shiftRegs_validIn_delay_186_0;
  reg                 shiftRegs_validIn_delay_187_0;
  reg                 shiftRegs_validIn_delay_188_0;
  reg                 shiftRegs_validIn_delay_189_0;
  reg                 shiftRegs_validIn_delay_190_0;
  reg                 shiftRegs_validIn_delay_191_0;
  reg                 shiftRegs_validIn_delay_192_0;
  reg                 shiftRegs_validIn_delay_193_0;
  reg                 shiftRegs_validIn_delay_194_0;
  reg                 shiftRegs_validIn_delay_195_0;
  reg                 shiftRegs_validIn_delay_196_0;
  reg                 shiftRegs_validIn_delay_197_0;
  reg                 shiftRegs_validIn_delay_198_0;
  reg                 shiftRegs_validIn_delay_199_0;
  reg                 shiftRegs_validIn_delay_200_0;
  reg                 shiftRegs_validIn_delay_201_0;
  reg                 shiftRegs_validIn_delay_202_0;
  reg                 shiftRegs_validIn_delay_203_0;
  reg                 shiftRegs_validIn_delay_204_0;
  reg                 shiftRegs_validIn_delay_205_0;
  reg                 shiftRegs_validIn_delay_206_0;
  reg                 shiftRegs_validIn_delay_207_0;
  reg                 shiftRegs_validIn_delay_208_0;
  reg                 shiftRegs_validIn_delay_209_0;
  reg                 shiftRegs_validIn_delay_210_0;
  reg                 shiftRegs_validIn_delay_211_0;
  reg                 shiftRegs_validIn_delay_212_0;
  reg                 shiftRegs_validIn_delay_213_0;
  reg                 shiftRegs_validIn_delay_214_0;
  reg                 shiftRegs_validIn_delay_215_0;
  reg                 shiftRegs_validIn_delay_216_0;
  reg                 shiftRegs_validIn_delay_217_0;
  reg                 shiftRegs_validIn_delay_218_0;
  reg                 shiftRegs_validIn_delay_219_0;
  reg                 shiftRegs_validIn_delay_220_0;
  reg                 shiftRegs_validIn_delay_221_0;
  reg                 shiftRegs_validIn_delay_222_0;
  reg                 shiftRegs_validIn_delay_223_0;
  reg                 shiftRegs_validIn_delay_224_0;
  reg                 shiftRegs_validIn_delay_225_0;
  reg                 shiftRegs_validIn_delay_226_0;
  reg                 shiftRegs_validIn_delay_227_0;
  reg                 shiftRegs_validIn_delay_228_0;
  reg                 shiftRegs_validIn_delay_229_0;
  reg                 shiftRegs_validIn_delay_230_0;
  reg                 shiftRegs_validIn_delay_231_0;
  reg                 shiftRegs_validIn_delay_232_0;
  reg                 shiftRegs_validIn_delay_233_0;
  reg                 shiftRegs_validIn_delay_234_0;
  reg                 shiftRegs_validIn_delay_235_0;
  reg                 shiftRegs_validIn_delay_236_0;
  reg                 shiftRegs_validIn_delay_237_0;
  reg                 shiftRegs_validIn_delay_238_0;
  reg                 shiftRegs_validIn_delay_239_0;
  reg                 shiftRegs_validIn_delay_240_0;
  reg                 shiftRegs_validIn_delay_241_0;
  reg                 shiftRegs_validIn_delay_242_0;
  reg                 shiftRegs_validIn_delay_243_0;
  reg                 shiftRegs_validIn_delay_244_0;
  reg                 shiftRegs_validIn_delay_245_0;
  reg                 shiftRegs_validIn_delay_246_0;
  reg                 shiftRegs_validIn_delay_247_0;
  reg                 shiftRegs_validIn_delay_248_0;
  reg                 shiftRegs_validIn_delay_249_0;
  reg                 shiftRegs_validIn_delay_250_0;
  reg                 shiftRegs_validIn_delay_251_0;
  reg                 shiftRegs_validIn_delay_252_0;
  reg                 shiftRegs_validIn_delay_253_0;
  reg                 shiftRegs_validIn_delay_254_0;
  reg                 shiftRegs_validOut_0;
  reg        [16:0]   shiftRegs_addressIn_delay_1_0;
  reg        [16:0]   shiftRegs_addressIn_delay_2_0;
  reg        [16:0]   shiftRegs_addressIn_delay_3_0;
  reg        [16:0]   shiftRegs_addressIn_delay_4_0;
  reg        [16:0]   shiftRegs_addressIn_delay_5_0;
  reg        [16:0]   shiftRegs_addressIn_delay_6_0;
  reg        [16:0]   shiftRegs_addressIn_delay_7_0;
  reg        [16:0]   shiftRegs_addressIn_delay_8_0;
  reg        [16:0]   shiftRegs_addressIn_delay_9_0;
  reg        [16:0]   shiftRegs_addressIn_delay_10_0;
  reg        [16:0]   shiftRegs_addressIn_delay_11_0;
  reg        [16:0]   shiftRegs_addressIn_delay_12_0;
  reg        [16:0]   shiftRegs_addressIn_delay_13_0;
  reg        [16:0]   shiftRegs_addressIn_delay_14_0;
  reg        [16:0]   shiftRegs_addressIn_delay_15_0;
  reg        [16:0]   shiftRegs_addressIn_delay_16_0;
  reg        [16:0]   shiftRegs_addressIn_delay_17_0;
  reg        [16:0]   shiftRegs_addressIn_delay_18_0;
  reg        [16:0]   shiftRegs_addressIn_delay_19_0;
  reg        [16:0]   shiftRegs_addressIn_delay_20_0;
  reg        [16:0]   shiftRegs_addressIn_delay_21_0;
  reg        [16:0]   shiftRegs_addressIn_delay_22_0;
  reg        [16:0]   shiftRegs_addressIn_delay_23_0;
  reg        [16:0]   shiftRegs_addressIn_delay_24_0;
  reg        [16:0]   shiftRegs_addressIn_delay_25_0;
  reg        [16:0]   shiftRegs_addressIn_delay_26_0;
  reg        [16:0]   shiftRegs_addressIn_delay_27_0;
  reg        [16:0]   shiftRegs_addressIn_delay_28_0;
  reg        [16:0]   shiftRegs_addressIn_delay_29_0;
  reg        [16:0]   shiftRegs_addressIn_delay_30_0;
  reg        [16:0]   shiftRegs_addressIn_delay_31_0;
  reg        [16:0]   shiftRegs_addressIn_delay_32_0;
  reg        [16:0]   shiftRegs_addressIn_delay_33_0;
  reg        [16:0]   shiftRegs_addressIn_delay_34_0;
  reg        [16:0]   shiftRegs_addressIn_delay_35_0;
  reg        [16:0]   shiftRegs_addressIn_delay_36_0;
  reg        [16:0]   shiftRegs_addressIn_delay_37_0;
  reg        [16:0]   shiftRegs_addressIn_delay_38_0;
  reg        [16:0]   shiftRegs_addressIn_delay_39_0;
  reg        [16:0]   shiftRegs_addressIn_delay_40_0;
  reg        [16:0]   shiftRegs_addressIn_delay_41_0;
  reg        [16:0]   shiftRegs_addressIn_delay_42_0;
  reg        [16:0]   shiftRegs_addressIn_delay_43_0;
  reg        [16:0]   shiftRegs_addressIn_delay_44_0;
  reg        [16:0]   shiftRegs_addressIn_delay_45_0;
  reg        [16:0]   shiftRegs_addressIn_delay_46_0;
  reg        [16:0]   shiftRegs_addressIn_delay_47_0;
  reg        [16:0]   shiftRegs_addressIn_delay_48_0;
  reg        [16:0]   shiftRegs_addressIn_delay_49_0;
  reg        [16:0]   shiftRegs_addressIn_delay_50_0;
  reg        [16:0]   shiftRegs_addressIn_delay_51_0;
  reg        [16:0]   shiftRegs_addressIn_delay_52_0;
  reg        [16:0]   shiftRegs_addressIn_delay_53_0;
  reg        [16:0]   shiftRegs_addressIn_delay_54_0;
  reg        [16:0]   shiftRegs_addressIn_delay_55_0;
  reg        [16:0]   shiftRegs_addressIn_delay_56_0;
  reg        [16:0]   shiftRegs_addressIn_delay_57_0;
  reg        [16:0]   shiftRegs_addressIn_delay_58_0;
  reg        [16:0]   shiftRegs_addressIn_delay_59_0;
  reg        [16:0]   shiftRegs_addressIn_delay_60_0;
  reg        [16:0]   shiftRegs_addressIn_delay_61_0;
  reg        [16:0]   shiftRegs_addressIn_delay_62_0;
  reg        [16:0]   shiftRegs_addressIn_delay_63_0;
  reg        [16:0]   shiftRegs_addressIn_delay_64_0;
  reg        [16:0]   shiftRegs_addressIn_delay_65_0;
  reg        [16:0]   shiftRegs_addressIn_delay_66_0;
  reg        [16:0]   shiftRegs_addressIn_delay_67_0;
  reg        [16:0]   shiftRegs_addressIn_delay_68_0;
  reg        [16:0]   shiftRegs_addressIn_delay_69_0;
  reg        [16:0]   shiftRegs_addressIn_delay_70_0;
  reg        [16:0]   shiftRegs_addressIn_delay_71_0;
  reg        [16:0]   shiftRegs_addressIn_delay_72_0;
  reg        [16:0]   shiftRegs_addressIn_delay_73_0;
  reg        [16:0]   shiftRegs_addressIn_delay_74_0;
  reg        [16:0]   shiftRegs_addressIn_delay_75_0;
  reg        [16:0]   shiftRegs_addressIn_delay_76_0;
  reg        [16:0]   shiftRegs_addressIn_delay_77_0;
  reg        [16:0]   shiftRegs_addressIn_delay_78_0;
  reg        [16:0]   shiftRegs_addressIn_delay_79_0;
  reg        [16:0]   shiftRegs_addressIn_delay_80_0;
  reg        [16:0]   shiftRegs_addressIn_delay_81_0;
  reg        [16:0]   shiftRegs_addressIn_delay_82_0;
  reg        [16:0]   shiftRegs_addressIn_delay_83_0;
  reg        [16:0]   shiftRegs_addressIn_delay_84_0;
  reg        [16:0]   shiftRegs_addressIn_delay_85_0;
  reg        [16:0]   shiftRegs_addressIn_delay_86_0;
  reg        [16:0]   shiftRegs_addressIn_delay_87_0;
  reg        [16:0]   shiftRegs_addressIn_delay_88_0;
  reg        [16:0]   shiftRegs_addressIn_delay_89_0;
  reg        [16:0]   shiftRegs_addressIn_delay_90_0;
  reg        [16:0]   shiftRegs_addressIn_delay_91_0;
  reg        [16:0]   shiftRegs_addressIn_delay_92_0;
  reg        [16:0]   shiftRegs_addressIn_delay_93_0;
  reg        [16:0]   shiftRegs_addressIn_delay_94_0;
  reg        [16:0]   shiftRegs_addressIn_delay_95_0;
  reg        [16:0]   shiftRegs_addressIn_delay_96_0;
  reg        [16:0]   shiftRegs_addressIn_delay_97_0;
  reg        [16:0]   shiftRegs_addressIn_delay_98_0;
  reg        [16:0]   shiftRegs_addressIn_delay_99_0;
  reg        [16:0]   shiftRegs_addressIn_delay_100_0;
  reg        [16:0]   shiftRegs_addressIn_delay_101_0;
  reg        [16:0]   shiftRegs_addressIn_delay_102_0;
  reg        [16:0]   shiftRegs_addressIn_delay_103_0;
  reg        [16:0]   shiftRegs_addressIn_delay_104_0;
  reg        [16:0]   shiftRegs_addressIn_delay_105_0;
  reg        [16:0]   shiftRegs_addressIn_delay_106_0;
  reg        [16:0]   shiftRegs_addressIn_delay_107_0;
  reg        [16:0]   shiftRegs_addressIn_delay_108_0;
  reg        [16:0]   shiftRegs_addressIn_delay_109_0;
  reg        [16:0]   shiftRegs_addressIn_delay_110_0;
  reg        [16:0]   shiftRegs_addressIn_delay_111_0;
  reg        [16:0]   shiftRegs_addressIn_delay_112_0;
  reg        [16:0]   shiftRegs_addressIn_delay_113_0;
  reg        [16:0]   shiftRegs_addressIn_delay_114_0;
  reg        [16:0]   shiftRegs_addressIn_delay_115_0;
  reg        [16:0]   shiftRegs_addressIn_delay_116_0;
  reg        [16:0]   shiftRegs_addressIn_delay_117_0;
  reg        [16:0]   shiftRegs_addressIn_delay_118_0;
  reg        [16:0]   shiftRegs_addressIn_delay_119_0;
  reg        [16:0]   shiftRegs_addressIn_delay_120_0;
  reg        [16:0]   shiftRegs_addressIn_delay_121_0;
  reg        [16:0]   shiftRegs_addressIn_delay_122_0;
  reg        [16:0]   shiftRegs_addressIn_delay_123_0;
  reg        [16:0]   shiftRegs_addressIn_delay_124_0;
  reg        [16:0]   shiftRegs_addressIn_delay_125_0;
  reg        [16:0]   shiftRegs_addressIn_delay_126_0;
  reg        [16:0]   shiftRegs_addressIn_delay_127_0;
  reg        [16:0]   shiftRegs_addressIn_delay_128_0;
  reg        [16:0]   shiftRegs_addressIn_delay_129_0;
  reg        [16:0]   shiftRegs_addressIn_delay_130_0;
  reg        [16:0]   shiftRegs_addressIn_delay_131_0;
  reg        [16:0]   shiftRegs_addressIn_delay_132_0;
  reg        [16:0]   shiftRegs_addressIn_delay_133_0;
  reg        [16:0]   shiftRegs_addressIn_delay_134_0;
  reg        [16:0]   shiftRegs_addressIn_delay_135_0;
  reg        [16:0]   shiftRegs_addressIn_delay_136_0;
  reg        [16:0]   shiftRegs_addressIn_delay_137_0;
  reg        [16:0]   shiftRegs_addressIn_delay_138_0;
  reg        [16:0]   shiftRegs_addressIn_delay_139_0;
  reg        [16:0]   shiftRegs_addressIn_delay_140_0;
  reg        [16:0]   shiftRegs_addressIn_delay_141_0;
  reg        [16:0]   shiftRegs_addressIn_delay_142_0;
  reg        [16:0]   shiftRegs_addressIn_delay_143_0;
  reg        [16:0]   shiftRegs_addressIn_delay_144_0;
  reg        [16:0]   shiftRegs_addressIn_delay_145_0;
  reg        [16:0]   shiftRegs_addressIn_delay_146_0;
  reg        [16:0]   shiftRegs_addressIn_delay_147_0;
  reg        [16:0]   shiftRegs_addressIn_delay_148_0;
  reg        [16:0]   shiftRegs_addressIn_delay_149_0;
  reg        [16:0]   shiftRegs_addressIn_delay_150_0;
  reg        [16:0]   shiftRegs_addressIn_delay_151_0;
  reg        [16:0]   shiftRegs_addressIn_delay_152_0;
  reg        [16:0]   shiftRegs_addressIn_delay_153_0;
  reg        [16:0]   shiftRegs_addressIn_delay_154_0;
  reg        [16:0]   shiftRegs_addressIn_delay_155_0;
  reg        [16:0]   shiftRegs_addressIn_delay_156_0;
  reg        [16:0]   shiftRegs_addressIn_delay_157_0;
  reg        [16:0]   shiftRegs_addressIn_delay_158_0;
  reg        [16:0]   shiftRegs_addressIn_delay_159_0;
  reg        [16:0]   shiftRegs_addressIn_delay_160_0;
  reg        [16:0]   shiftRegs_addressIn_delay_161_0;
  reg        [16:0]   shiftRegs_addressIn_delay_162_0;
  reg        [16:0]   shiftRegs_addressIn_delay_163_0;
  reg        [16:0]   shiftRegs_addressIn_delay_164_0;
  reg        [16:0]   shiftRegs_addressIn_delay_165_0;
  reg        [16:0]   shiftRegs_addressIn_delay_166_0;
  reg        [16:0]   shiftRegs_addressIn_delay_167_0;
  reg        [16:0]   shiftRegs_addressIn_delay_168_0;
  reg        [16:0]   shiftRegs_addressIn_delay_169_0;
  reg        [16:0]   shiftRegs_addressIn_delay_170_0;
  reg        [16:0]   shiftRegs_addressIn_delay_171_0;
  reg        [16:0]   shiftRegs_addressIn_delay_172_0;
  reg        [16:0]   shiftRegs_addressIn_delay_173_0;
  reg        [16:0]   shiftRegs_addressIn_delay_174_0;
  reg        [16:0]   shiftRegs_addressIn_delay_175_0;
  reg        [16:0]   shiftRegs_addressIn_delay_176_0;
  reg        [16:0]   shiftRegs_addressIn_delay_177_0;
  reg        [16:0]   shiftRegs_addressIn_delay_178_0;
  reg        [16:0]   shiftRegs_addressIn_delay_179_0;
  reg        [16:0]   shiftRegs_addressIn_delay_180_0;
  reg        [16:0]   shiftRegs_addressIn_delay_181_0;
  reg        [16:0]   shiftRegs_addressIn_delay_182_0;
  reg        [16:0]   shiftRegs_addressIn_delay_183_0;
  reg        [16:0]   shiftRegs_addressIn_delay_184_0;
  reg        [16:0]   shiftRegs_addressIn_delay_185_0;
  reg        [16:0]   shiftRegs_addressIn_delay_186_0;
  reg        [16:0]   shiftRegs_addressIn_delay_187_0;
  reg        [16:0]   shiftRegs_addressIn_delay_188_0;
  reg        [16:0]   shiftRegs_addressIn_delay_189_0;
  reg        [16:0]   shiftRegs_addressIn_delay_190_0;
  reg        [16:0]   shiftRegs_addressIn_delay_191_0;
  reg        [16:0]   shiftRegs_addressIn_delay_192_0;
  reg        [16:0]   shiftRegs_addressIn_delay_193_0;
  reg        [16:0]   shiftRegs_addressIn_delay_194_0;
  reg        [16:0]   shiftRegs_addressIn_delay_195_0;
  reg        [16:0]   shiftRegs_addressIn_delay_196_0;
  reg        [16:0]   shiftRegs_addressIn_delay_197_0;
  reg        [16:0]   shiftRegs_addressIn_delay_198_0;
  reg        [16:0]   shiftRegs_addressIn_delay_199_0;
  reg        [16:0]   shiftRegs_addressIn_delay_200_0;
  reg        [16:0]   shiftRegs_addressIn_delay_201_0;
  reg        [16:0]   shiftRegs_addressIn_delay_202_0;
  reg        [16:0]   shiftRegs_addressIn_delay_203_0;
  reg        [16:0]   shiftRegs_addressIn_delay_204_0;
  reg        [16:0]   shiftRegs_addressIn_delay_205_0;
  reg        [16:0]   shiftRegs_addressIn_delay_206_0;
  reg        [16:0]   shiftRegs_addressIn_delay_207_0;
  reg        [16:0]   shiftRegs_addressIn_delay_208_0;
  reg        [16:0]   shiftRegs_addressIn_delay_209_0;
  reg        [16:0]   shiftRegs_addressIn_delay_210_0;
  reg        [16:0]   shiftRegs_addressIn_delay_211_0;
  reg        [16:0]   shiftRegs_addressIn_delay_212_0;
  reg        [16:0]   shiftRegs_addressIn_delay_213_0;
  reg        [16:0]   shiftRegs_addressIn_delay_214_0;
  reg        [16:0]   shiftRegs_addressIn_delay_215_0;
  reg        [16:0]   shiftRegs_addressIn_delay_216_0;
  reg        [16:0]   shiftRegs_addressIn_delay_217_0;
  reg        [16:0]   shiftRegs_addressIn_delay_218_0;
  reg        [16:0]   shiftRegs_addressIn_delay_219_0;
  reg        [16:0]   shiftRegs_addressIn_delay_220_0;
  reg        [16:0]   shiftRegs_addressIn_delay_221_0;
  reg        [16:0]   shiftRegs_addressIn_delay_222_0;
  reg        [16:0]   shiftRegs_addressIn_delay_223_0;
  reg        [16:0]   shiftRegs_addressIn_delay_224_0;
  reg        [16:0]   shiftRegs_addressIn_delay_225_0;
  reg        [16:0]   shiftRegs_addressIn_delay_226_0;
  reg        [16:0]   shiftRegs_addressIn_delay_227_0;
  reg        [16:0]   shiftRegs_addressIn_delay_228_0;
  reg        [16:0]   shiftRegs_addressIn_delay_229_0;
  reg        [16:0]   shiftRegs_addressIn_delay_230_0;
  reg        [16:0]   shiftRegs_addressIn_delay_231_0;
  reg        [16:0]   shiftRegs_addressIn_delay_232_0;
  reg        [16:0]   shiftRegs_addressIn_delay_233_0;
  reg        [16:0]   shiftRegs_addressIn_delay_234_0;
  reg        [16:0]   shiftRegs_addressIn_delay_235_0;
  reg        [16:0]   shiftRegs_addressIn_delay_236_0;
  reg        [16:0]   shiftRegs_addressIn_delay_237_0;
  reg        [16:0]   shiftRegs_addressIn_delay_238_0;
  reg        [16:0]   shiftRegs_addressIn_delay_239_0;
  reg        [16:0]   shiftRegs_addressIn_delay_240_0;
  reg        [16:0]   shiftRegs_addressIn_delay_241_0;
  reg        [16:0]   shiftRegs_addressIn_delay_242_0;
  reg        [16:0]   shiftRegs_addressIn_delay_243_0;
  reg        [16:0]   shiftRegs_addressIn_delay_244_0;
  reg        [16:0]   shiftRegs_addressIn_delay_245_0;
  reg        [16:0]   shiftRegs_addressIn_delay_246_0;
  reg        [16:0]   shiftRegs_addressIn_delay_247_0;
  reg        [16:0]   shiftRegs_addressIn_delay_248_0;
  reg        [16:0]   shiftRegs_addressIn_delay_249_0;
  reg        [16:0]   shiftRegs_addressIn_delay_250_0;
  reg        [16:0]   shiftRegs_addressIn_delay_251_0;
  reg        [16:0]   shiftRegs_addressIn_delay_252_0;
  reg        [16:0]   shiftRegs_addressIn_delay_253_0;
  reg        [16:0]   shiftRegs_addressIn_delay_254_0;
  reg        [16:0]   shiftRegs_addressOut_0;
  reg                 shiftRegs_validOut_delay_1_0;
  reg                 shiftRegs_validOut_delay_2_0;
  reg                 shiftRegs_validOut_delay_3_0;
  reg                 shiftRegs_validOut_delay_4_0;
  reg                 shiftRegs_validOutFull_0;
  reg        [16:0]   shiftRegs_addressOut_delay_1_0;
  reg        [16:0]   shiftRegs_addressOut_delay_2_0;
  reg        [16:0]   shiftRegs_addressOut_delay_3_0;
  reg        [16:0]   shiftRegs_addressOut_delay_4_0;
  reg        [16:0]   shiftRegs_addressOutFull_0;
  reg                 outputValid;
  reg        [376:0]  pAddPort_0_s_regNext_X;
  reg        [376:0]  pAddPort_0_s_regNext_Y;
  reg        [376:0]  pAddPort_0_s_regNext_Z;
  reg        [376:0]  pAddPort_0_s_regNext_T;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg                 flushing_flushCnt_willIncrement;
  wire                flushing_flushCnt_willClear;
  reg        [16:0]   flushing_flushCnt_valueNext;
  reg        [16:0]   flushing_flushCnt_value;
  reg                 flushing_flushCnt_willOverflowIfInc;
  wire                flushing_flushCnt_willOverflow;
  reg                 stage1_NCnt_willIncrement;
  reg                 stage1_NCnt_willClear;
  reg        [31:0]   stage1_NCnt_valueNext;
  reg        [31:0]   stage1_NCnt_value;
  reg                 stage1_NCnt_willOverflowIfInc;
  wire                stage1_NCnt_willOverflow;
  reg                 stage1_GCnt_willIncrement;
  wire                stage1_GCnt_willClear;
  reg        [4:0]    stage1_GCnt_valueNext;
  reg        [4:0]    stage1_GCnt_value;
  reg                 stage1_GCnt_willOverflowIfInc;
  wire                stage1_GCnt_willOverflow;
  reg                 stage1_waitReg;
  reg                 stage1_emptyCnt_willIncrement;
  reg                 stage1_emptyCnt_willClear;
  reg        [8:0]    stage1_emptyCnt_valueNext;
  reg        [8:0]    stage1_emptyCnt_value;
  reg                 stage1_emptyCnt_willOverflowIfInc;
  wire                stage1_emptyCnt_willOverflow;
  reg                 stage1_needAdd1_0;
  wire       [13:0]   stage1_inputBarrelID_0;
  wire       [12:0]   _zz_stage1_inputBarrelIDAbs_0;
  wire       [11:0]   stage1_inputBarrelIDAbs_0;
  reg                 _zz_stage1_inputValid_0;
  reg                 _zz_stage1_inputValid_0_1;
  reg                 _zz_stage1_inputValid_0_2;
  reg                 _zz_stage1_inputValid_0_3;
  reg                 _zz_stage1_inputValid_0_4;
  reg                 stage1_inputValid_0;
  reg        [16:0]   _zz_stage1_inputAddress_0;
  reg        [16:0]   _zz_stage1_inputAddress_0_1;
  reg        [16:0]   _zz_stage1_inputAddress_0_2;
  reg        [16:0]   _zz_stage1_inputAddress_0_3;
  reg        [16:0]   _zz_stage1_inputAddress_0_4;
  reg        [16:0]   stage1_inputAddress_0;
  reg                 _zz_stage1_inputData_0_X;
  reg                 _zz_stage1_inputData_0_X_1;
  reg                 _zz_stage1_inputData_0_X_2;
  reg                 _zz_stage1_inputData_0_X_3;
  reg                 _zz_stage1_inputData_0_X_4;
  reg                 _zz_stage1_inputData_0_X_5;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_1_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_2_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_3_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_4_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_5_T;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_X;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z;
  reg        [376:0]  dataInBuffer_bufferOut_payload_fragment_P_delay_6_T;
  wire       [376:0]  stage1_inputData_0_X;
  wire       [376:0]  stage1_inputData_0_Y;
  wire       [376:0]  stage1_inputData_0_Z;
  wire       [376:0]  stage1_inputData_0_T;
  reg                 stage2_wCnt_willDecrement;
  wire                stage2_wCnt_willClear;
  reg        [11:0]   stage2_wCnt_valueNext;
  reg        [11:0]   stage2_wCnt_value;
  reg                 stage2_wCnt_willUnderflowIfDec;
  wire                stage2_wCnt_willUnderflow;
  reg                 stage2_GCnt_willIncrement;
  wire                stage2_GCnt_willClear;
  reg        [4:0]    stage2_GCnt_valueNext;
  reg        [4:0]    stage2_GCnt_value;
  reg                 stage2_GCnt_willOverflowIfInc;
  wire                stage2_GCnt_willOverflow;
  reg                 stage2_calCnt_willDecrement;
  wire                stage2_calCnt_willClear;
  reg        [1:0]    stage2_calCnt_valueNext;
  reg        [1:0]    stage2_calCnt_value;
  reg                 stage2_calCnt_willUnderflowIfDec;
  wire                stage2_calCnt_willUnderflow;
  reg                 stage2_waitReg;
  reg                 stage2_waitCnt_willIncrement;
  wire                stage2_waitCnt_willClear;
  reg        [8:0]    stage2_waitCnt_valueNext;
  reg        [8:0]    stage2_waitCnt_value;
  reg                 stage2_waitCnt_willOverflowIfInc;
  wire                stage2_waitCnt_willOverflow;
  reg                 stage3_GCnt_willDecrement;
  wire                stage3_GCnt_willClear;
  reg        [4:0]    stage3_GCnt_valueNext;
  reg        [4:0]    stage3_GCnt_value;
  reg                 stage3_GCnt_willUnderflowIfDec;
  wire                stage3_GCnt_willUnderflow;
  reg                 stage3_doubleCnt_willIncrement;
  wire                stage3_doubleCnt_willClear;
  reg        [3:0]    stage3_doubleCnt_valueNext;
  reg        [3:0]    stage3_doubleCnt_value;
  reg                 stage3_doubleCnt_willOverflowIfInc;
  wire                stage3_doubleCnt_willOverflow;
  reg                 stage3_doubleWaitCnt_willIncrement;
  wire                stage3_doubleWaitCnt_willClear;
  reg        [8:0]    stage3_doubleWaitCnt_valueNext;
  reg        [8:0]    stage3_doubleWaitCnt_value;
  reg                 stage3_doubleWaitCnt_willOverflowIfInc;
  wire                stage3_doubleWaitCnt_willOverflow;
  reg                 stage3_addReg;
  reg                 stage3_addWaitCnt_willIncrement;
  wire                stage3_addWaitCnt_willClear;
  reg        [8:0]    stage3_addWaitCnt_valueNext;
  reg        [8:0]    stage3_addWaitCnt_value;
  reg                 stage3_addWaitCnt_willOverflowIfInc;
  wire                stage3_addWaitCnt_willOverflow;
  reg        [3:0]    fsm_stateReg;
  reg        [3:0]    fsm_stateNext;
  reg                 stage1_inputValid_0_delay_1;
  reg                 stage1_inputValid_0_delay_2;
  reg                 stage1_inputValid_0_delay_3;
  reg                 stage1_inputValid_0_delay_4;
  reg                 stage1_inputValid_0_delay_5;
  reg        [16:0]   stage1_inputAddress_0_delay_1;
  reg        [16:0]   stage1_inputAddress_0_delay_2;
  reg        [16:0]   stage1_inputAddress_0_delay_3;
  reg        [16:0]   stage1_inputAddress_0_delay_4;
  reg        [16:0]   stage1_inputAddress_0_delay_5;
  reg        [376:0]  stage1_inputData_0_delay_1_X;
  reg        [376:0]  stage1_inputData_0_delay_1_Y;
  reg        [376:0]  stage1_inputData_0_delay_1_Z;
  reg        [376:0]  stage1_inputData_0_delay_1_T;
  reg        [376:0]  stage1_inputData_0_delay_2_X;
  reg        [376:0]  stage1_inputData_0_delay_2_Y;
  reg        [376:0]  stage1_inputData_0_delay_2_Z;
  reg        [376:0]  stage1_inputData_0_delay_2_T;
  reg        [376:0]  stage1_inputData_0_delay_3_X;
  reg        [376:0]  stage1_inputData_0_delay_3_Y;
  reg        [376:0]  stage1_inputData_0_delay_3_Z;
  reg        [376:0]  stage1_inputData_0_delay_3_T;
  reg        [376:0]  stage1_inputData_0_delay_4_X;
  reg        [376:0]  stage1_inputData_0_delay_4_Y;
  reg        [376:0]  stage1_inputData_0_delay_4_Z;
  reg        [376:0]  stage1_inputData_0_delay_4_T;
  reg        [376:0]  stage1_inputData_0_delay_5_X;
  reg        [376:0]  stage1_inputData_0_delay_5_Y;
  reg        [376:0]  stage1_inputData_0_delay_5_Z;
  reg        [376:0]  stage1_inputData_0_delay_5_T;
  reg                 _zz_io_dataIn_0_valid;
  reg                 _zz_io_dataIn_0_valid_1;
  reg                 _zz_io_dataIn_0_valid_2;
  reg                 _zz_io_dataIn_0_valid_3;
  reg                 _zz_io_dataIn_0_valid_4;
  reg                 _zz_io_dataIn_0_valid_5;
  reg                 _zz_io_dataIn_0_valid_6;
  reg                 _zz_io_dataIn_0_valid_7;
  reg                 _zz_io_dataIn_0_valid_8;
  reg                 _zz_io_dataIn_0_valid_9;
  reg                 _zz_io_dataIn_0_valid_10;
  reg                 _zz_io_dataIn_0_valid_11;
  reg                 _zz_io_dataIn_0_valid_12;
  reg                 _zz_io_dataIn_0_valid_13;
  reg                 _zz_io_dataIn_0_valid_14;
  reg                 _zz_io_dataIn_0_valid_15;
  reg                 _zz_io_dataIn_0_valid_16;
  reg                 _zz_io_dataIn_0_valid_17;
  reg                 _zz_io_dataIn_0_valid_18;
  reg                 _zz_io_dataIn_0_valid_19;
  reg                 _zz_io_dataIn_0_valid_20;
  reg                 _zz_io_dataIn_0_valid_21;
  reg                 _zz_io_dataIn_0_valid_22;
  reg                 _zz_io_dataIn_0_valid_23;
  reg                 _zz_io_dataIn_0_valid_24;
  reg                 _zz_io_dataIn_0_valid_25;
  reg                 _zz_io_dataIn_0_valid_26;
  reg                 _zz_io_dataIn_0_valid_27;
  reg                 _zz_io_dataIn_0_valid_28;
  reg                 _zz_io_dataIn_0_valid_29;
  reg                 _zz_io_dataIn_0_valid_30;
  reg                 _zz_io_dataIn_0_valid_31;
  reg                 _zz_io_dataIn_0_valid_32;
  reg                 _zz_io_dataIn_0_valid_33;
  reg                 _zz_io_dataIn_0_valid_34;
  reg                 _zz_io_dataIn_0_payload_a_X;
  reg                 _zz_io_dataIn_0_payload_a_X_1;
  reg                 _zz_io_dataIn_0_payload_a_X_2;
  reg                 _zz_io_dataIn_0_payload_a_X_3;
  reg                 _zz_io_dataIn_0_payload_a_X_4;
  reg                 _zz_io_dataIn_0_payload_a_X_5;
  reg                 _zz_io_dataIn_0_payload_a_X_6;
  reg                 _zz_io_dataIn_0_payload_a_X_7;
  reg                 _zz_io_dataIn_0_payload_a_X_8;
  reg                 _zz_io_dataIn_0_payload_a_X_9;
  reg                 _zz_io_dataIn_0_payload_a_X_10;
  reg                 _zz_io_dataIn_0_payload_a_X_11;
  reg                 _zz_io_dataIn_0_payload_a_X_12;
  reg                 _zz_io_dataIn_0_payload_a_X_13;
  reg                 _zz_io_dataIn_0_payload_a_X_14;
  reg                 _zz_io_dataIn_0_payload_a_X_15;
  reg                 _zz_io_dataIn_0_payload_a_X_16;
  reg                 _zz_io_dataIn_0_payload_a_X_17;
  reg                 _zz_io_dataIn_0_payload_a_X_18;
  reg                 _zz_io_dataIn_0_payload_a_X_19;
  reg                 _zz_io_dataIn_0_payload_a_X_20;
  reg                 _zz_io_dataIn_0_payload_a_X_21;
  reg                 _zz_io_dataIn_0_payload_a_X_22;
  reg                 _zz_io_dataIn_0_payload_a_X_23;
  reg                 _zz_io_dataIn_0_payload_a_X_24;
  reg                 _zz_io_dataIn_0_payload_a_X_25;
  reg                 _zz_io_dataIn_0_payload_a_X_26;
  reg                 _zz_io_dataIn_0_payload_a_X_27;
  reg                 _zz_io_dataIn_0_payload_a_X_28;
  reg                 _zz_io_dataIn_0_payload_a_X_29;
  reg                 _zz_io_dataIn_0_payload_a_X_30;
  reg                 _zz_io_dataIn_0_payload_a_X_31;
  reg                 _zz_io_dataIn_0_payload_a_X_32;
  reg                 _zz_io_dataIn_0_payload_a_X_33;
  reg                 _zz_io_dataIn_0_payload_a_X_34;
  reg        [376:0]  stage1_inputData_0_delay_1_X_1;
  reg        [376:0]  stage1_inputData_0_delay_1_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_1_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_1_T_1;
  reg        [376:0]  stage1_inputData_0_delay_2_X_1;
  reg        [376:0]  stage1_inputData_0_delay_2_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_2_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_2_T_1;
  reg        [376:0]  stage1_inputData_0_delay_3_X_1;
  reg        [376:0]  stage1_inputData_0_delay_3_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_3_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_3_T_1;
  reg        [376:0]  stage1_inputData_0_delay_4_X_1;
  reg        [376:0]  stage1_inputData_0_delay_4_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_4_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_4_T_1;
  reg        [376:0]  stage1_inputData_0_delay_5_X_1;
  reg        [376:0]  stage1_inputData_0_delay_5_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_5_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_5_T_1;
  reg        [376:0]  stage1_inputData_0_delay_6_X;
  reg        [376:0]  stage1_inputData_0_delay_6_Y;
  reg        [376:0]  stage1_inputData_0_delay_6_Z;
  reg        [376:0]  stage1_inputData_0_delay_6_T;
  reg        [376:0]  stage1_inputData_0_delay_7_X;
  reg        [376:0]  stage1_inputData_0_delay_7_Y;
  reg        [376:0]  stage1_inputData_0_delay_7_Z;
  reg        [376:0]  stage1_inputData_0_delay_7_T;
  reg        [376:0]  stage1_inputData_0_delay_8_X;
  reg        [376:0]  stage1_inputData_0_delay_8_Y;
  reg        [376:0]  stage1_inputData_0_delay_8_Z;
  reg        [376:0]  stage1_inputData_0_delay_8_T;
  reg        [376:0]  stage1_inputData_0_delay_9_X;
  reg        [376:0]  stage1_inputData_0_delay_9_Y;
  reg        [376:0]  stage1_inputData_0_delay_9_Z;
  reg        [376:0]  stage1_inputData_0_delay_9_T;
  reg        [376:0]  stage1_inputData_0_delay_10_X;
  reg        [376:0]  stage1_inputData_0_delay_10_Y;
  reg        [376:0]  stage1_inputData_0_delay_10_Z;
  reg        [376:0]  stage1_inputData_0_delay_10_T;
  reg        [376:0]  stage1_inputData_0_delay_11_X;
  reg        [376:0]  stage1_inputData_0_delay_11_Y;
  reg        [376:0]  stage1_inputData_0_delay_11_Z;
  reg        [376:0]  stage1_inputData_0_delay_11_T;
  reg        [376:0]  stage1_inputData_0_delay_12_X;
  reg        [376:0]  stage1_inputData_0_delay_12_Y;
  reg        [376:0]  stage1_inputData_0_delay_12_Z;
  reg        [376:0]  stage1_inputData_0_delay_12_T;
  reg        [376:0]  stage1_inputData_0_delay_13_X;
  reg        [376:0]  stage1_inputData_0_delay_13_Y;
  reg        [376:0]  stage1_inputData_0_delay_13_Z;
  reg        [376:0]  stage1_inputData_0_delay_13_T;
  reg        [376:0]  stage1_inputData_0_delay_14_X;
  reg        [376:0]  stage1_inputData_0_delay_14_Y;
  reg        [376:0]  stage1_inputData_0_delay_14_Z;
  reg        [376:0]  stage1_inputData_0_delay_14_T;
  reg        [376:0]  stage1_inputData_0_delay_15_X;
  reg        [376:0]  stage1_inputData_0_delay_15_Y;
  reg        [376:0]  stage1_inputData_0_delay_15_Z;
  reg        [376:0]  stage1_inputData_0_delay_15_T;
  reg        [376:0]  stage1_inputData_0_delay_16_X;
  reg        [376:0]  stage1_inputData_0_delay_16_Y;
  reg        [376:0]  stage1_inputData_0_delay_16_Z;
  reg        [376:0]  stage1_inputData_0_delay_16_T;
  reg        [376:0]  stage1_inputData_0_delay_17_X;
  reg        [376:0]  stage1_inputData_0_delay_17_Y;
  reg        [376:0]  stage1_inputData_0_delay_17_Z;
  reg        [376:0]  stage1_inputData_0_delay_17_T;
  reg        [376:0]  stage1_inputData_0_delay_18_X;
  reg        [376:0]  stage1_inputData_0_delay_18_Y;
  reg        [376:0]  stage1_inputData_0_delay_18_Z;
  reg        [376:0]  stage1_inputData_0_delay_18_T;
  reg        [376:0]  stage1_inputData_0_delay_19_X;
  reg        [376:0]  stage1_inputData_0_delay_19_Y;
  reg        [376:0]  stage1_inputData_0_delay_19_Z;
  reg        [376:0]  stage1_inputData_0_delay_19_T;
  reg        [376:0]  stage1_inputData_0_delay_20_X;
  reg        [376:0]  stage1_inputData_0_delay_20_Y;
  reg        [376:0]  stage1_inputData_0_delay_20_Z;
  reg        [376:0]  stage1_inputData_0_delay_20_T;
  reg        [376:0]  stage1_inputData_0_delay_21_X;
  reg        [376:0]  stage1_inputData_0_delay_21_Y;
  reg        [376:0]  stage1_inputData_0_delay_21_Z;
  reg        [376:0]  stage1_inputData_0_delay_21_T;
  reg        [376:0]  stage1_inputData_0_delay_22_X;
  reg        [376:0]  stage1_inputData_0_delay_22_Y;
  reg        [376:0]  stage1_inputData_0_delay_22_Z;
  reg        [376:0]  stage1_inputData_0_delay_22_T;
  reg        [376:0]  stage1_inputData_0_delay_23_X;
  reg        [376:0]  stage1_inputData_0_delay_23_Y;
  reg        [376:0]  stage1_inputData_0_delay_23_Z;
  reg        [376:0]  stage1_inputData_0_delay_23_T;
  reg        [376:0]  stage1_inputData_0_delay_24_X;
  reg        [376:0]  stage1_inputData_0_delay_24_Y;
  reg        [376:0]  stage1_inputData_0_delay_24_Z;
  reg        [376:0]  stage1_inputData_0_delay_24_T;
  reg        [376:0]  stage1_inputData_0_delay_25_X;
  reg        [376:0]  stage1_inputData_0_delay_25_Y;
  reg        [376:0]  stage1_inputData_0_delay_25_Z;
  reg        [376:0]  stage1_inputData_0_delay_25_T;
  reg        [376:0]  stage1_inputData_0_delay_26_X;
  reg        [376:0]  stage1_inputData_0_delay_26_Y;
  reg        [376:0]  stage1_inputData_0_delay_26_Z;
  reg        [376:0]  stage1_inputData_0_delay_26_T;
  reg        [376:0]  stage1_inputData_0_delay_27_X;
  reg        [376:0]  stage1_inputData_0_delay_27_Y;
  reg        [376:0]  stage1_inputData_0_delay_27_Z;
  reg        [376:0]  stage1_inputData_0_delay_27_T;
  reg        [376:0]  stage1_inputData_0_delay_28_X;
  reg        [376:0]  stage1_inputData_0_delay_28_Y;
  reg        [376:0]  stage1_inputData_0_delay_28_Z;
  reg        [376:0]  stage1_inputData_0_delay_28_T;
  reg        [376:0]  stage1_inputData_0_delay_29_X;
  reg        [376:0]  stage1_inputData_0_delay_29_Y;
  reg        [376:0]  stage1_inputData_0_delay_29_Z;
  reg        [376:0]  stage1_inputData_0_delay_29_T;
  reg        [376:0]  stage1_inputData_0_delay_30_X;
  reg        [376:0]  stage1_inputData_0_delay_30_Y;
  reg        [376:0]  stage1_inputData_0_delay_30_Z;
  reg        [376:0]  stage1_inputData_0_delay_30_T;
  reg        [376:0]  stage1_inputData_0_delay_31_X;
  reg        [376:0]  stage1_inputData_0_delay_31_Y;
  reg        [376:0]  stage1_inputData_0_delay_31_Z;
  reg        [376:0]  stage1_inputData_0_delay_31_T;
  reg        [376:0]  stage1_inputData_0_delay_32_X;
  reg        [376:0]  stage1_inputData_0_delay_32_Y;
  reg        [376:0]  stage1_inputData_0_delay_32_Z;
  reg        [376:0]  stage1_inputData_0_delay_32_T;
  reg        [376:0]  stage1_inputData_0_delay_33_X;
  reg        [376:0]  stage1_inputData_0_delay_33_Y;
  reg        [376:0]  stage1_inputData_0_delay_33_Z;
  reg        [376:0]  stage1_inputData_0_delay_33_T;
  reg        [376:0]  stage1_inputData_0_delay_34_X;
  reg        [376:0]  stage1_inputData_0_delay_34_Y;
  reg        [376:0]  stage1_inputData_0_delay_34_Z;
  reg        [376:0]  stage1_inputData_0_delay_34_T;
  reg        [376:0]  stage1_inputData_0_delay_35_X;
  reg        [376:0]  stage1_inputData_0_delay_35_Y;
  reg        [376:0]  stage1_inputData_0_delay_35_Z;
  reg        [376:0]  stage1_inputData_0_delay_35_T;
  reg        [376:0]  pAddPort_0_s_delay_1_X;
  reg        [376:0]  pAddPort_0_s_delay_1_Y;
  reg        [376:0]  pAddPort_0_s_delay_1_Z;
  reg        [376:0]  pAddPort_0_s_delay_1_T;
  reg        [376:0]  pAddPort_0_s_delay_2_X;
  reg        [376:0]  pAddPort_0_s_delay_2_Y;
  reg        [376:0]  pAddPort_0_s_delay_2_Z;
  reg        [376:0]  pAddPort_0_s_delay_2_T;
  reg        [376:0]  pAddPort_0_s_delay_3_X;
  reg        [376:0]  pAddPort_0_s_delay_3_Y;
  reg        [376:0]  pAddPort_0_s_delay_3_Z;
  reg        [376:0]  pAddPort_0_s_delay_3_T;
  reg        [376:0]  pAddPort_0_s_delay_4_X;
  reg        [376:0]  pAddPort_0_s_delay_4_Y;
  reg        [376:0]  pAddPort_0_s_delay_4_Z;
  reg        [376:0]  pAddPort_0_s_delay_4_T;
  reg        [376:0]  pAddPort_0_s_delay_5_X;
  reg        [376:0]  pAddPort_0_s_delay_5_Y;
  reg        [376:0]  pAddPort_0_s_delay_5_Z;
  reg        [376:0]  pAddPort_0_s_delay_5_T;
  reg        [376:0]  pAddPort_0_s_delay_6_X;
  reg        [376:0]  pAddPort_0_s_delay_6_Y;
  reg        [376:0]  pAddPort_0_s_delay_6_Z;
  reg        [376:0]  pAddPort_0_s_delay_6_T;
  reg        [376:0]  pAddPort_0_s_delay_7_X;
  reg        [376:0]  pAddPort_0_s_delay_7_Y;
  reg        [376:0]  pAddPort_0_s_delay_7_Z;
  reg        [376:0]  pAddPort_0_s_delay_7_T;
  reg        [376:0]  pAddPort_0_s_delay_8_X;
  reg        [376:0]  pAddPort_0_s_delay_8_Y;
  reg        [376:0]  pAddPort_0_s_delay_8_Z;
  reg        [376:0]  pAddPort_0_s_delay_8_T;
  reg        [376:0]  pAddPort_0_s_delay_9_X;
  reg        [376:0]  pAddPort_0_s_delay_9_Y;
  reg        [376:0]  pAddPort_0_s_delay_9_Z;
  reg        [376:0]  pAddPort_0_s_delay_9_T;
  reg        [376:0]  pAddPort_0_s_delay_10_X;
  reg        [376:0]  pAddPort_0_s_delay_10_Y;
  reg        [376:0]  pAddPort_0_s_delay_10_Z;
  reg        [376:0]  pAddPort_0_s_delay_10_T;
  reg        [376:0]  pAddPort_0_s_delay_11_X;
  reg        [376:0]  pAddPort_0_s_delay_11_Y;
  reg        [376:0]  pAddPort_0_s_delay_11_Z;
  reg        [376:0]  pAddPort_0_s_delay_11_T;
  reg        [376:0]  pAddPort_0_s_delay_12_X;
  reg        [376:0]  pAddPort_0_s_delay_12_Y;
  reg        [376:0]  pAddPort_0_s_delay_12_Z;
  reg        [376:0]  pAddPort_0_s_delay_12_T;
  reg        [376:0]  pAddPort_0_s_delay_13_X;
  reg        [376:0]  pAddPort_0_s_delay_13_Y;
  reg        [376:0]  pAddPort_0_s_delay_13_Z;
  reg        [376:0]  pAddPort_0_s_delay_13_T;
  reg        [376:0]  pAddPort_0_s_delay_14_X;
  reg        [376:0]  pAddPort_0_s_delay_14_Y;
  reg        [376:0]  pAddPort_0_s_delay_14_Z;
  reg        [376:0]  pAddPort_0_s_delay_14_T;
  reg        [376:0]  pAddPort_0_s_delay_15_X;
  reg        [376:0]  pAddPort_0_s_delay_15_Y;
  reg        [376:0]  pAddPort_0_s_delay_15_Z;
  reg        [376:0]  pAddPort_0_s_delay_15_T;
  reg        [376:0]  pAddPort_0_s_delay_16_X;
  reg        [376:0]  pAddPort_0_s_delay_16_Y;
  reg        [376:0]  pAddPort_0_s_delay_16_Z;
  reg        [376:0]  pAddPort_0_s_delay_16_T;
  reg        [376:0]  pAddPort_0_s_delay_17_X;
  reg        [376:0]  pAddPort_0_s_delay_17_Y;
  reg        [376:0]  pAddPort_0_s_delay_17_Z;
  reg        [376:0]  pAddPort_0_s_delay_17_T;
  reg        [376:0]  pAddPort_0_s_delay_18_X;
  reg        [376:0]  pAddPort_0_s_delay_18_Y;
  reg        [376:0]  pAddPort_0_s_delay_18_Z;
  reg        [376:0]  pAddPort_0_s_delay_18_T;
  reg        [376:0]  pAddPort_0_s_delay_19_X;
  reg        [376:0]  pAddPort_0_s_delay_19_Y;
  reg        [376:0]  pAddPort_0_s_delay_19_Z;
  reg        [376:0]  pAddPort_0_s_delay_19_T;
  reg        [376:0]  pAddPort_0_s_delay_20_X;
  reg        [376:0]  pAddPort_0_s_delay_20_Y;
  reg        [376:0]  pAddPort_0_s_delay_20_Z;
  reg        [376:0]  pAddPort_0_s_delay_20_T;
  reg        [376:0]  pAddPort_0_s_delay_21_X;
  reg        [376:0]  pAddPort_0_s_delay_21_Y;
  reg        [376:0]  pAddPort_0_s_delay_21_Z;
  reg        [376:0]  pAddPort_0_s_delay_21_T;
  reg        [376:0]  pAddPort_0_s_delay_22_X;
  reg        [376:0]  pAddPort_0_s_delay_22_Y;
  reg        [376:0]  pAddPort_0_s_delay_22_Z;
  reg        [376:0]  pAddPort_0_s_delay_22_T;
  reg        [376:0]  pAddPort_0_s_delay_23_X;
  reg        [376:0]  pAddPort_0_s_delay_23_Y;
  reg        [376:0]  pAddPort_0_s_delay_23_Z;
  reg        [376:0]  pAddPort_0_s_delay_23_T;
  reg        [376:0]  pAddPort_0_s_delay_24_X;
  reg        [376:0]  pAddPort_0_s_delay_24_Y;
  reg        [376:0]  pAddPort_0_s_delay_24_Z;
  reg        [376:0]  pAddPort_0_s_delay_24_T;
  reg        [376:0]  pAddPort_0_s_delay_25_X;
  reg        [376:0]  pAddPort_0_s_delay_25_Y;
  reg        [376:0]  pAddPort_0_s_delay_25_Z;
  reg        [376:0]  pAddPort_0_s_delay_25_T;
  reg        [376:0]  pAddPort_0_s_delay_26_X;
  reg        [376:0]  pAddPort_0_s_delay_26_Y;
  reg        [376:0]  pAddPort_0_s_delay_26_Z;
  reg        [376:0]  pAddPort_0_s_delay_26_T;
  reg        [376:0]  pAddPort_0_s_delay_27_X;
  reg        [376:0]  pAddPort_0_s_delay_27_Y;
  reg        [376:0]  pAddPort_0_s_delay_27_Z;
  reg        [376:0]  pAddPort_0_s_delay_27_T;
  reg        [376:0]  pAddPort_0_s_delay_28_X;
  reg        [376:0]  pAddPort_0_s_delay_28_Y;
  reg        [376:0]  pAddPort_0_s_delay_28_Z;
  reg        [376:0]  pAddPort_0_s_delay_28_T;
  reg        [376:0]  pAddPort_0_s_delay_29_X;
  reg        [376:0]  pAddPort_0_s_delay_29_Y;
  reg        [376:0]  pAddPort_0_s_delay_29_Z;
  reg        [376:0]  pAddPort_0_s_delay_29_T;
  reg        [376:0]  pAddPort_0_s_delay_30_X;
  reg        [376:0]  pAddPort_0_s_delay_30_Y;
  reg        [376:0]  pAddPort_0_s_delay_30_Z;
  reg        [376:0]  pAddPort_0_s_delay_30_T;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_1;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_2;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_3;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_4;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_5;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_6;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_7;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_8;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_9;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_10;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_11;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_12;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_13;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_14;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_15;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_16;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_17;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_18;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_19;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_20;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_21;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_22;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_23;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_24;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_25;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_26;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_27;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_28;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_29;
  reg        [16:0]   shiftRegs_addressOutFull_0_delay_30;
  reg                 _zz_io_dataIn_1_valid;
  reg                 _zz_io_dataIn_1_valid_1;
  reg                 _zz_io_dataIn_1_valid_2;
  reg                 _zz_io_dataIn_1_valid_3;
  reg                 _zz_io_dataIn_1_valid_4;
  reg                 _zz_io_dataIn_1_valid_5;
  reg                 _zz_io_dataIn_1_valid_6;
  reg                 _zz_io_dataIn_1_valid_7;
  reg                 _zz_io_dataIn_1_valid_8;
  reg                 _zz_io_dataIn_1_valid_9;
  reg                 _zz_io_dataIn_1_valid_10;
  reg                 _zz_io_dataIn_1_valid_11;
  reg                 _zz_io_dataIn_1_valid_12;
  reg                 _zz_io_dataIn_1_valid_13;
  reg                 _zz_io_dataIn_1_valid_14;
  reg                 _zz_io_dataIn_1_valid_15;
  reg                 _zz_io_dataIn_1_valid_16;
  reg                 _zz_io_dataIn_1_valid_17;
  reg                 _zz_io_dataIn_1_valid_18;
  reg                 _zz_io_dataIn_1_valid_19;
  reg                 _zz_io_dataIn_1_valid_20;
  reg                 _zz_io_dataIn_1_valid_21;
  reg                 _zz_io_dataIn_1_valid_22;
  reg                 _zz_io_dataIn_1_valid_23;
  reg                 _zz_io_dataIn_1_valid_24;
  reg                 _zz_io_dataIn_1_valid_25;
  reg                 _zz_io_dataIn_1_valid_26;
  reg                 _zz_io_dataIn_1_valid_27;
  reg                 _zz_io_dataIn_1_valid_28;
  reg                 _zz_io_dataIn_1_valid_29;
  reg                 _zz_io_dataIn_1_valid_30;
  reg                 _zz_io_dataIn_1_valid_31;
  reg                 _zz_io_dataIn_1_valid_32;
  reg                 _zz_io_dataIn_1_valid_33;
  reg                 _zz_io_dataIn_1_valid_34;
  reg        [376:0]  stage1_inputData_0_delay_1_X_2;
  reg        [376:0]  stage1_inputData_0_delay_1_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_1_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_1_T_2;
  reg        [376:0]  stage1_inputData_0_delay_2_X_2;
  reg        [376:0]  stage1_inputData_0_delay_2_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_2_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_2_T_2;
  reg        [376:0]  stage1_inputData_0_delay_3_X_2;
  reg        [376:0]  stage1_inputData_0_delay_3_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_3_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_3_T_2;
  reg        [376:0]  stage1_inputData_0_delay_4_X_2;
  reg        [376:0]  stage1_inputData_0_delay_4_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_4_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_4_T_2;
  reg        [376:0]  stage1_inputData_0_delay_5_X_2;
  reg        [376:0]  stage1_inputData_0_delay_5_Y_2;
  reg        [376:0]  stage1_inputData_0_delay_5_Z_2;
  reg        [376:0]  stage1_inputData_0_delay_5_T_2;
  reg        [376:0]  stage1_inputData_0_delay_6_X_1;
  reg        [376:0]  stage1_inputData_0_delay_6_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_6_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_6_T_1;
  reg        [376:0]  stage1_inputData_0_delay_7_X_1;
  reg        [376:0]  stage1_inputData_0_delay_7_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_7_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_7_T_1;
  reg        [376:0]  stage1_inputData_0_delay_8_X_1;
  reg        [376:0]  stage1_inputData_0_delay_8_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_8_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_8_T_1;
  reg        [376:0]  stage1_inputData_0_delay_9_X_1;
  reg        [376:0]  stage1_inputData_0_delay_9_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_9_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_9_T_1;
  reg        [376:0]  stage1_inputData_0_delay_10_X_1;
  reg        [376:0]  stage1_inputData_0_delay_10_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_10_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_10_T_1;
  reg        [376:0]  stage1_inputData_0_delay_11_X_1;
  reg        [376:0]  stage1_inputData_0_delay_11_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_11_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_11_T_1;
  reg        [376:0]  stage1_inputData_0_delay_12_X_1;
  reg        [376:0]  stage1_inputData_0_delay_12_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_12_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_12_T_1;
  reg        [376:0]  stage1_inputData_0_delay_13_X_1;
  reg        [376:0]  stage1_inputData_0_delay_13_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_13_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_13_T_1;
  reg        [376:0]  stage1_inputData_0_delay_14_X_1;
  reg        [376:0]  stage1_inputData_0_delay_14_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_14_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_14_T_1;
  reg        [376:0]  stage1_inputData_0_delay_15_X_1;
  reg        [376:0]  stage1_inputData_0_delay_15_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_15_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_15_T_1;
  reg        [376:0]  stage1_inputData_0_delay_16_X_1;
  reg        [376:0]  stage1_inputData_0_delay_16_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_16_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_16_T_1;
  reg        [376:0]  stage1_inputData_0_delay_17_X_1;
  reg        [376:0]  stage1_inputData_0_delay_17_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_17_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_17_T_1;
  reg        [376:0]  stage1_inputData_0_delay_18_X_1;
  reg        [376:0]  stage1_inputData_0_delay_18_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_18_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_18_T_1;
  reg        [376:0]  stage1_inputData_0_delay_19_X_1;
  reg        [376:0]  stage1_inputData_0_delay_19_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_19_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_19_T_1;
  reg        [376:0]  stage1_inputData_0_delay_20_X_1;
  reg        [376:0]  stage1_inputData_0_delay_20_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_20_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_20_T_1;
  reg        [376:0]  stage1_inputData_0_delay_21_X_1;
  reg        [376:0]  stage1_inputData_0_delay_21_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_21_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_21_T_1;
  reg        [376:0]  stage1_inputData_0_delay_22_X_1;
  reg        [376:0]  stage1_inputData_0_delay_22_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_22_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_22_T_1;
  reg        [376:0]  stage1_inputData_0_delay_23_X_1;
  reg        [376:0]  stage1_inputData_0_delay_23_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_23_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_23_T_1;
  reg        [376:0]  stage1_inputData_0_delay_24_X_1;
  reg        [376:0]  stage1_inputData_0_delay_24_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_24_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_24_T_1;
  reg        [376:0]  stage1_inputData_0_delay_25_X_1;
  reg        [376:0]  stage1_inputData_0_delay_25_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_25_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_25_T_1;
  reg        [376:0]  stage1_inputData_0_delay_26_X_1;
  reg        [376:0]  stage1_inputData_0_delay_26_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_26_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_26_T_1;
  reg        [376:0]  stage1_inputData_0_delay_27_X_1;
  reg        [376:0]  stage1_inputData_0_delay_27_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_27_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_27_T_1;
  reg        [376:0]  stage1_inputData_0_delay_28_X_1;
  reg        [376:0]  stage1_inputData_0_delay_28_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_28_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_28_T_1;
  reg        [376:0]  stage1_inputData_0_delay_29_X_1;
  reg        [376:0]  stage1_inputData_0_delay_29_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_29_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_29_T_1;
  reg        [376:0]  stage1_inputData_0_delay_30_X_1;
  reg        [376:0]  stage1_inputData_0_delay_30_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_30_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_30_T_1;
  reg        [376:0]  stage1_inputData_0_delay_31_X_1;
  reg        [376:0]  stage1_inputData_0_delay_31_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_31_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_31_T_1;
  reg        [376:0]  stage1_inputData_0_delay_32_X_1;
  reg        [376:0]  stage1_inputData_0_delay_32_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_32_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_32_T_1;
  reg        [376:0]  stage1_inputData_0_delay_33_X_1;
  reg        [376:0]  stage1_inputData_0_delay_33_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_33_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_33_T_1;
  reg        [376:0]  stage1_inputData_0_delay_34_X_1;
  reg        [376:0]  stage1_inputData_0_delay_34_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_34_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_34_T_1;
  reg        [376:0]  stage1_inputData_0_delay_35_X_1;
  reg        [376:0]  stage1_inputData_0_delay_35_Y_1;
  reg        [376:0]  stage1_inputData_0_delay_35_Z_1;
  reg        [376:0]  stage1_inputData_0_delay_35_T_1;
  reg        [16:0]   stage1_inputAddress_0_delay_1_1;
  reg        [16:0]   stage1_inputAddress_0_delay_2_1;
  reg        [16:0]   stage1_inputAddress_0_delay_3_1;
  reg        [16:0]   stage1_inputAddress_0_delay_4_1;
  reg        [16:0]   stage1_inputAddress_0_delay_5_1;
  reg        [16:0]   stage1_inputAddress_0_delay_6;
  reg        [16:0]   stage1_inputAddress_0_delay_7;
  reg        [16:0]   stage1_inputAddress_0_delay_8;
  reg        [16:0]   stage1_inputAddress_0_delay_9;
  reg        [16:0]   stage1_inputAddress_0_delay_10;
  reg        [16:0]   stage1_inputAddress_0_delay_11;
  reg        [16:0]   stage1_inputAddress_0_delay_12;
  reg        [16:0]   stage1_inputAddress_0_delay_13;
  reg        [16:0]   stage1_inputAddress_0_delay_14;
  reg        [16:0]   stage1_inputAddress_0_delay_15;
  reg        [16:0]   stage1_inputAddress_0_delay_16;
  reg        [16:0]   stage1_inputAddress_0_delay_17;
  reg        [16:0]   stage1_inputAddress_0_delay_18;
  reg        [16:0]   stage1_inputAddress_0_delay_19;
  reg        [16:0]   stage1_inputAddress_0_delay_20;
  reg        [16:0]   stage1_inputAddress_0_delay_21;
  reg        [16:0]   stage1_inputAddress_0_delay_22;
  reg        [16:0]   stage1_inputAddress_0_delay_23;
  reg        [16:0]   stage1_inputAddress_0_delay_24;
  reg        [16:0]   stage1_inputAddress_0_delay_25;
  reg        [16:0]   stage1_inputAddress_0_delay_26;
  reg        [16:0]   stage1_inputAddress_0_delay_27;
  reg        [16:0]   stage1_inputAddress_0_delay_28;
  reg        [16:0]   stage1_inputAddress_0_delay_29;
  reg        [16:0]   stage1_inputAddress_0_delay_30;
  reg        [16:0]   stage1_inputAddress_0_delay_31;
  reg        [16:0]   stage1_inputAddress_0_delay_32;
  reg        [16:0]   stage1_inputAddress_0_delay_33;
  reg        [16:0]   stage1_inputAddress_0_delay_34;
  reg        [16:0]   stage1_inputAddress_0_delay_35;
  wire                when_Pippenger_l153;
  wire                when_Pippenger_l168;
  reg                 _zz_io_state_1;
  reg                 _zz_io_state_1_1;
  reg                 _zz_io_state_1_2;
  reg                 _zz_io_state_1_3;
  reg                 _zz_io_state_1_4;
  reg                 _zz_io_state_1_5;
  reg                 _zz_io_state_1_6;
  reg                 _zz_io_state_1_7;
  reg                 _zz_io_state_1_8;
  reg                 _zz_io_state_1_9;
  reg                 _zz_io_state_1_10;
  reg                 _zz_io_state_1_11;
  reg                 _zz_io_state_1_12;
  reg                 _zz_io_state_1_13;
  reg                 _zz_io_state_1_14;
  reg                 _zz_io_state_1_15;
  reg                 _zz_io_state_1_16;
  reg                 _zz_io_state_1_17;
  reg                 _zz_io_state_1_18;
  reg                 _zz_io_state_1_19;
  reg                 _zz_io_state_1_20;
  reg                 _zz_io_state_1_21;
  reg                 _zz_io_state_1_22;
  reg                 _zz_io_state_1_23;
  reg                 _zz_io_state_1_24;
  reg                 _zz_io_state_1_25;
  reg                 _zz_io_state_1_26;
  reg                 _zz_io_state_1_27;
  reg                 _zz_io_state_1_28;
  reg                 _zz_io_state_1_29;
  reg                 _zz_io_state_1_30;
  reg                 _zz_io_state_1_31;
  reg                 _zz_io_state_1_32;
  reg                 _zz_io_state_1_33;
  reg                 _zz_io_state_1_34;
  reg                 _zz_io_state_1_35;
  reg                 _zz_io_state_1_36;
  reg                 _zz_io_state_1_37;
  reg                 _zz_io_state_1_38;
  reg                 _zz_io_dataIn_1_valid_35;
  reg                 _zz_io_dataIn_1_valid_36;
  reg                 _zz_io_dataIn_1_valid_37;
  reg                 _zz_io_dataIn_1_valid_38;
  reg                 _zz_io_dataIn_1_valid_39;
  reg                 _zz_io_dataIn_1_valid_40;
  reg                 _zz_io_dataIn_1_valid_41;
  reg                 _zz_io_dataIn_1_valid_42;
  reg                 _zz_io_dataIn_1_valid_43;
  reg                 _zz_io_dataIn_1_valid_44;
  reg                 _zz_io_dataIn_1_valid_45;
  reg                 _zz_io_dataIn_1_valid_46;
  reg                 _zz_io_dataIn_1_valid_47;
  reg                 _zz_io_dataIn_1_valid_48;
  reg                 _zz_io_dataIn_1_valid_49;
  reg                 _zz_io_dataIn_1_valid_50;
  reg                 _zz_io_dataIn_1_valid_51;
  reg                 _zz_io_dataIn_1_valid_52;
  reg                 _zz_io_dataIn_1_valid_53;
  reg                 _zz_io_dataIn_1_valid_54;
  reg                 _zz_io_dataIn_1_valid_55;
  reg                 _zz_io_dataIn_1_valid_56;
  reg                 _zz_io_dataIn_1_valid_57;
  reg                 _zz_io_dataIn_1_valid_58;
  reg                 _zz_io_dataIn_1_valid_59;
  reg                 _zz_io_dataIn_1_valid_60;
  reg                 _zz_io_dataIn_1_valid_61;
  reg                 _zz_io_dataIn_1_valid_62;
  reg                 _zz_io_dataIn_1_valid_63;
  reg                 _zz_io_dataIn_1_valid_64;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_X;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_Y;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_Z;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_T;
  reg        [16:0]   _zz_io_dataIn_1_payload_address;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_1;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_2;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_3;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_4;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_5;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_6;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_7;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_8;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_9;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_10;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_11;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_12;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_13;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_14;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_15;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_16;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_17;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_18;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_19;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_20;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_21;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_22;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_23;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_24;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_25;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_26;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_27;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_28;
  reg        [16:0]   _zz_io_dataIn_1_payload_address_29;
  wire                when_Pippenger_l207;
  reg                 _zz_io_dataIn_1_valid_65;
  reg                 _zz_io_dataIn_1_valid_66;
  reg                 _zz_io_dataIn_1_valid_67;
  reg                 _zz_io_dataIn_1_valid_68;
  reg                 _zz_io_dataIn_1_valid_69;
  reg                 _zz_io_dataIn_1_valid_70;
  reg                 _zz_io_dataIn_1_valid_71;
  reg                 _zz_io_dataIn_1_valid_72;
  reg                 _zz_io_dataIn_1_valid_73;
  reg                 _zz_io_dataIn_1_valid_74;
  reg                 _zz_io_dataIn_1_valid_75;
  reg                 _zz_io_dataIn_1_valid_76;
  reg                 _zz_io_dataIn_1_valid_77;
  reg                 _zz_io_dataIn_1_valid_78;
  reg                 _zz_io_dataIn_1_valid_79;
  reg                 _zz_io_dataIn_1_valid_80;
  reg                 _zz_io_dataIn_1_valid_81;
  reg                 _zz_io_dataIn_1_valid_82;
  reg                 _zz_io_dataIn_1_valid_83;
  reg                 _zz_io_dataIn_1_valid_84;
  reg                 _zz_io_dataIn_1_valid_85;
  reg                 _zz_io_dataIn_1_valid_86;
  reg                 _zz_io_dataIn_1_valid_87;
  reg                 _zz_io_dataIn_1_valid_88;
  reg                 _zz_io_dataIn_1_valid_89;
  reg                 _zz_io_dataIn_1_valid_90;
  reg                 _zz_io_dataIn_1_valid_91;
  reg                 _zz_io_dataIn_1_valid_92;
  reg                 _zz_io_dataIn_1_valid_93;
  reg                 _zz_io_dataIn_1_valid_94;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_X_1;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_Y_1;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_Z_1;
  reg        [376:0]  pippenger_1_dataRam_0_io_rData_1_regNext_T_1;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_30;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_31;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_32;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_33;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_34;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_35;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_36;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_37;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_38;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_39;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_40;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_41;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_42;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_43;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_44;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_45;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_46;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_47;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_48;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_49;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_50;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_51;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_52;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_53;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_54;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_55;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_56;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_57;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_58;
  reg        [4:0]    _zz_io_dataIn_1_payload_address_59;
  wire                when_Pippenger_l249;
  `ifndef SYNTHESIS
  reg [63:0] fsm_stateReg_string;
  reg [63:0] fsm_stateNext_string;
  `endif


  assign _zz_dataInBuffer_dataReg_fragment_K = (dataInBuffer_dataReg_fragment_K >>> 13);
  assign _zz_flushing_flushCnt_valueNext_1 = flushing_flushCnt_willIncrement;
  assign _zz_flushing_flushCnt_valueNext = {16'd0, _zz_flushing_flushCnt_valueNext_1};
  assign _zz_stage1_NCnt_valueNext_1 = stage1_NCnt_willIncrement;
  assign _zz_stage1_NCnt_valueNext = {31'd0, _zz_stage1_NCnt_valueNext_1};
  assign _zz_stage1_GCnt_valueNext_1 = stage1_GCnt_willIncrement;
  assign _zz_stage1_GCnt_valueNext = {4'd0, _zz_stage1_GCnt_valueNext_1};
  assign _zz_stage1_emptyCnt_valueNext_1 = stage1_emptyCnt_willIncrement;
  assign _zz_stage1_emptyCnt_valueNext = {8'd0, _zz_stage1_emptyCnt_valueNext_1};
  assign _zz_stage1_inputBarrelID_0 = dataInBuffer_bufferOut_payload_fragment_K[12:0];
  assign _zz_stage1_inputBarrelID_0_2 = {1'b0,stage1_needAdd1_0};
  assign _zz_stage1_inputBarrelID_0_1 = {12'd0, _zz_stage1_inputBarrelID_0_2};
  assign _zz__zz_stage1_inputBarrelIDAbs_0 = stage1_inputBarrelID_0[12:0];
  assign _zz_stage1_inputBarrelIDAbs_0_1 = (_zz_stage1_inputBarrelIDAbs_0_2 + _zz_stage1_inputBarrelIDAbs_0_4);
  assign _zz_stage1_inputBarrelIDAbs_0_2 = (_zz_stage1_inputBarrelIDAbs_0[12] ? _zz_stage1_inputBarrelIDAbs_0_3 : _zz_stage1_inputBarrelIDAbs_0);
  assign _zz_stage1_inputBarrelIDAbs_0_3 = (~ _zz_stage1_inputBarrelIDAbs_0);
  assign _zz_stage1_inputBarrelIDAbs_0_5 = _zz_stage1_inputBarrelIDAbs_0[12];
  assign _zz_stage1_inputBarrelIDAbs_0_4 = {12'd0, _zz_stage1_inputBarrelIDAbs_0_5};
  assign _zz__zz_stage1_inputValid_0 = stage1_inputBarrelID_0[12:0];
  assign _zz_stage2_wCnt_valueNext_1 = stage2_wCnt_willDecrement;
  assign _zz_stage2_wCnt_valueNext = {11'd0, _zz_stage2_wCnt_valueNext_1};
  assign _zz_stage2_GCnt_valueNext_1 = stage2_GCnt_willIncrement;
  assign _zz_stage2_GCnt_valueNext = {4'd0, _zz_stage2_GCnt_valueNext_1};
  assign _zz_stage2_calCnt_valueNext_1 = stage2_calCnt_willDecrement;
  assign _zz_stage2_calCnt_valueNext = {1'd0, _zz_stage2_calCnt_valueNext_1};
  assign _zz_stage2_waitCnt_valueNext_1 = stage2_waitCnt_willIncrement;
  assign _zz_stage2_waitCnt_valueNext = {8'd0, _zz_stage2_waitCnt_valueNext_1};
  assign _zz_stage3_GCnt_valueNext_1 = stage3_GCnt_willDecrement;
  assign _zz_stage3_GCnt_valueNext = {4'd0, _zz_stage3_GCnt_valueNext_1};
  assign _zz_stage3_doubleCnt_valueNext_1 = stage3_doubleCnt_willIncrement;
  assign _zz_stage3_doubleCnt_valueNext = {3'd0, _zz_stage3_doubleCnt_valueNext_1};
  assign _zz_stage3_doubleWaitCnt_valueNext_1 = stage3_doubleWaitCnt_willIncrement;
  assign _zz_stage3_doubleWaitCnt_valueNext = {8'd0, _zz_stage3_doubleWaitCnt_valueNext_1};
  assign _zz_stage3_addWaitCnt_valueNext_1 = stage3_addWaitCnt_willIncrement;
  assign _zz_stage3_addWaitCnt_valueNext = {8'd0, _zz_stage3_addWaitCnt_valueNext_1};
  assign _zz_io_address_0_1 = (stage2_wCnt_value + _zz_io_address_0_2);
  assign _zz_io_address_0 = _zz_io_address_0_1;
  assign _zz_io_address_0_2 = {10'd0, stage2_calCnt_value};
  assign _zz_io_address_1_1 = (stage2_wCnt_value + _zz_io_address_1_2);
  assign _zz_io_address_1 = _zz_io_address_1_1;
  assign _zz_io_address_1_2 = {10'd0, stage2_calCnt_value};
  assign _zz__zz_io_dataIn_1_payload_address_1 = (stage2_wCnt_value + _zz__zz_io_dataIn_1_payload_address_2);
  assign _zz__zz_io_dataIn_1_payload_address = _zz__zz_io_dataIn_1_payload_address_1;
  assign _zz__zz_io_dataIn_1_payload_address_2 = {10'd0, stage2_calCnt_value};
  assign _zz_io_address_1_3 = (stage3_GCnt_value - _zz_io_address_1_4);
  assign _zz_io_address_1_5 = stage3_addWaitCnt_value[0];
  assign _zz_io_address_1_4 = {4'd0, _zz_io_address_1_5};
  assign _zz__zz_io_dataIn_1_payload_address_30_1 = stage3_addWaitCnt_value[0];
  assign _zz__zz_io_dataIn_1_payload_address_30 = {4'd0, _zz__zz_io_dataIn_1_payload_address_30_1};
  StateRam stateRam_0 (
    .io_we_0      (stateRam_0_io_we_0           ), //i
    .io_we_1      (stateRam_0_io_we_1           ), //i
    .io_address_0 (stateRam_0_io_address_0[16:0]), //i
    .io_address_1 (stateRam_0_io_address_1[16:0]), //i
    .io_state_0   (stateRam_0_io_state_0        ), //o
    .io_state_1   (stateRam_0_io_state_1        ), //o
    .io_flush     (stateRam_0_io_flush          ), //i
    .io_flushCnt  (stateRam_0_io_flushCnt[16:0] ), //i
    .clk          (clk                          ), //i
    .resetn       (resetn                       )  //i
  );
  DataRam dataRam_0 (
    .io_we_0      (dataRam_0_io_we_0            ), //i
    .io_we_1      (dataRam_0_io_we_1            ), //i
    .io_address_0 (dataRam_0_io_address_0[16:0] ), //i
    .io_address_1 (dataRam_0_io_address_1[16:0] ), //i
    .io_wData_0_X (dataRam_0_io_wData_0_X[376:0]), //i
    .io_wData_0_Y (dataRam_0_io_wData_0_Y[376:0]), //i
    .io_wData_0_Z (dataRam_0_io_wData_0_Z[376:0]), //i
    .io_wData_0_T (dataRam_0_io_wData_0_T[376:0]), //i
    .io_wData_1_X (dataRam_0_io_wData_1_X[376:0]), //i
    .io_wData_1_Y (dataRam_0_io_wData_1_Y[376:0]), //i
    .io_wData_1_Z (dataRam_0_io_wData_1_Z[376:0]), //i
    .io_wData_1_T (dataRam_0_io_wData_1_T[376:0]), //i
    .io_state_0   (1'b1                         ), //i
    .io_state_1   (dataRam_0_io_state_1         ), //i
    .io_rData_0_X (dataRam_0_io_rData_0_X[376:0]), //o
    .io_rData_0_Y (dataRam_0_io_rData_0_Y[376:0]), //o
    .io_rData_0_Z (dataRam_0_io_rData_0_Z[376:0]), //o
    .io_rData_0_T (dataRam_0_io_rData_0_T[376:0]), //o
    .io_rData_1_X (dataRam_0_io_rData_1_X[376:0]), //o
    .io_rData_1_Y (dataRam_0_io_rData_1_Y[376:0]), //o
    .io_rData_1_Z (dataRam_0_io_rData_1_Z[376:0]), //o
    .io_rData_1_T (dataRam_0_io_rData_1_T[376:0]), //o
    .io_pInit_X   (io_pInit_X[376:0]            ), //i
    .io_pInit_Y   (io_pInit_Y[376:0]            ), //i
    .io_pInit_Z   (io_pInit_Z[376:0]            ), //i
    .io_pInit_T   (io_pInit_T[376:0]            ), //i
    .clk          (clk                          ), //i
    .resetn       (resetn                       )  //i
  );
  DWSRFIFO fifo_0 (
    .io_dataIn_0_valid           (fifo_0_io_dataIn_0_valid                ), //i
    .io_dataIn_0_payload_a_X     (fifo_0_io_dataIn_0_payload_a_X[376:0]   ), //i
    .io_dataIn_0_payload_a_Y     (fifo_0_io_dataIn_0_payload_a_Y[376:0]   ), //i
    .io_dataIn_0_payload_a_Z     (fifo_0_io_dataIn_0_payload_a_Z[376:0]   ), //i
    .io_dataIn_0_payload_a_T     (fifo_0_io_dataIn_0_payload_a_T[376:0]   ), //i
    .io_dataIn_0_payload_b_X     (fifo_0_io_dataIn_0_payload_b_X[376:0]   ), //i
    .io_dataIn_0_payload_b_Y     (fifo_0_io_dataIn_0_payload_b_Y[376:0]   ), //i
    .io_dataIn_0_payload_b_Z     (fifo_0_io_dataIn_0_payload_b_Z[376:0]   ), //i
    .io_dataIn_0_payload_b_T     (fifo_0_io_dataIn_0_payload_b_T[376:0]   ), //i
    .io_dataIn_0_payload_address (fifo_0_io_dataIn_0_payload_address[16:0]), //i
    .io_dataIn_1_valid           (fifo_0_io_dataIn_1_valid                ), //i
    .io_dataIn_1_payload_a_X     (fifo_0_io_dataIn_1_payload_a_X[376:0]   ), //i
    .io_dataIn_1_payload_a_Y     (fifo_0_io_dataIn_1_payload_a_Y[376:0]   ), //i
    .io_dataIn_1_payload_a_Z     (fifo_0_io_dataIn_1_payload_a_Z[376:0]   ), //i
    .io_dataIn_1_payload_a_T     (fifo_0_io_dataIn_1_payload_a_T[376:0]   ), //i
    .io_dataIn_1_payload_b_X     (fifo_0_io_dataIn_1_payload_b_X[376:0]   ), //i
    .io_dataIn_1_payload_b_Y     (fifo_0_io_dataIn_1_payload_b_Y[376:0]   ), //i
    .io_dataIn_1_payload_b_Z     (fifo_0_io_dataIn_1_payload_b_Z[376:0]   ), //i
    .io_dataIn_1_payload_b_T     (fifo_0_io_dataIn_1_payload_b_T[376:0]   ), //i
    .io_dataIn_1_payload_address (fifo_0_io_dataIn_1_payload_address[16:0]), //i
    .io_dataOut_valid            (fifo_0_io_dataOut_valid                 ), //o
    .io_dataOut_payload_a_X      (fifo_0_io_dataOut_payload_a_X[376:0]    ), //o
    .io_dataOut_payload_a_Y      (fifo_0_io_dataOut_payload_a_Y[376:0]    ), //o
    .io_dataOut_payload_a_Z      (fifo_0_io_dataOut_payload_a_Z[376:0]    ), //o
    .io_dataOut_payload_a_T      (fifo_0_io_dataOut_payload_a_T[376:0]    ), //o
    .io_dataOut_payload_b_X      (fifo_0_io_dataOut_payload_b_X[376:0]    ), //o
    .io_dataOut_payload_b_Y      (fifo_0_io_dataOut_payload_b_Y[376:0]    ), //o
    .io_dataOut_payload_b_Z      (fifo_0_io_dataOut_payload_b_Z[376:0]    ), //o
    .io_dataOut_payload_b_T      (fifo_0_io_dataOut_payload_b_T[376:0]    ), //o
    .io_dataOut_payload_address  (fifo_0_io_dataOut_payload_address[16:0] ), //o
    .clk                         (clk                                     ), //i
    .resetn                      (resetn                                  )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_flushing : fsm_stateReg_string = "flushing";
      fsm_enumDef_stage1 : fsm_stateReg_string = "stage1  ";
      fsm_enumDef_stage2 : fsm_stateReg_string = "stage2  ";
      fsm_enumDef_stage3 : fsm_stateReg_string = "stage3  ";
      default : fsm_stateReg_string = "????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_flushing : fsm_stateNext_string = "flushing";
      fsm_enumDef_stage1 : fsm_stateNext_string = "stage1  ";
      fsm_enumDef_stage2 : fsm_stateNext_string = "stage2  ";
      fsm_enumDef_stage3 : fsm_stateNext_string = "stage3  ";
      default : fsm_stateNext_string = "????????";
    endcase
  end
  `endif

  assign dataInBuffer_bufferOut_valid = dataInBuffer_validReg;
  assign dataInBuffer_bufferOut_payload_last = dataInBuffer_dataReg_last;
  assign dataInBuffer_bufferOut_payload_fragment_P_X = dataInBuffer_dataReg_fragment_P_X;
  assign dataInBuffer_bufferOut_payload_fragment_P_Y = dataInBuffer_dataReg_fragment_P_Y;
  assign dataInBuffer_bufferOut_payload_fragment_P_Z = dataInBuffer_dataReg_fragment_P_Z;
  assign dataInBuffer_bufferOut_payload_fragment_P_T = dataInBuffer_dataReg_fragment_P_T;
  assign dataInBuffer_bufferOut_payload_fragment_K = dataInBuffer_dataReg_fragment_K;
  assign io_dataIn_ready = ((! dataInBuffer_validReg) || dataInBuffer_bufferOut_ready);
  always @(*) begin
    dataInBuffer_bufferOut_ready = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          if(dataInBuffer_bufferOut_valid) begin
            if(stage1_GCnt_willOverflowIfInc) begin
              dataInBuffer_bufferOut_ready = 1'b1;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataInBuffer_shift = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          dataInBuffer_shift = 1'b1;
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_we_0 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_0_io_we_0 = shiftRegs_validOut_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_we_1 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_0_io_we_1 = stage1_inputValid_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_address_0 = 17'bxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_0_io_address_0 = shiftRegs_addressOut_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_0_io_address_0 = {stage2_GCnt_value,_zz_io_address_0};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_address_1 = 17'bxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        stateRam_0_io_address_1 = stage1_inputAddress_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_flush = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_0_io_flush = stage2_calCnt_willUnderflowIfDec;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
        stateRam_0_io_flush = 1'b1;
      end
    endcase
  end

  always @(*) begin
    stateRam_0_io_flushCnt = 17'bxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        stateRam_0_io_flushCnt = {stage2_GCnt_value,stage2_wCnt_value};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
        stateRam_0_io_flushCnt = flushing_flushCnt_value;
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_we_0 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_we_0 = ((! stateRam_0_io_state_0) && shiftRegs_validOutFull_0);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_we_0 = shiftRegs_validOutFull_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_we_0 = shiftRegs_validOutFull_0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_we_1 = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_we_1 = ((! stateRam_0_io_state_1) && stage1_inputValid_0_delay_5);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_address_0 = 17'bxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_address_0 = shiftRegs_addressOutFull_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_address_0 = shiftRegs_addressOutFull_0;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_address_0 = shiftRegs_addressOutFull_0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_address_1 = 17'bxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_address_1 = stage1_inputAddress_0_delay_5;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_address_1 = {stage2_GCnt_value,_zz_io_address_1};
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_address_1 = {_zz_io_address_1_3,12'h001};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_0_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_0_X = pAddPort_0_s_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_wData_0_X = pAddPort_0_s_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_wData_0_X = pAddPort_0_s_X;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_0_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_0_Y = pAddPort_0_s_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_wData_0_Y = pAddPort_0_s_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_wData_0_Y = pAddPort_0_s_Y;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_0_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_0_Z = pAddPort_0_s_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_wData_0_Z = pAddPort_0_s_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_wData_0_Z = pAddPort_0_s_Z;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_0_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_0_T = pAddPort_0_s_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_wData_0_T = pAddPort_0_s_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        dataRam_0_io_wData_0_T = pAddPort_0_s_T;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_1_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_1_X = stage1_inputData_0_delay_5_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_1_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_1_Y = stage1_inputData_0_delay_5_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_1_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_1_Z = stage1_inputData_0_delay_5_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_wData_1_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        dataRam_0_io_wData_1_T = stage1_inputData_0_delay_5_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    dataRam_0_io_state_1 = 1'b1;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        dataRam_0_io_state_1 = _zz_io_state_1_38;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_valid = _zz_io_dataIn_0_valid_34;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_a_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_a_X = (_zz_io_dataIn_0_payload_a_X_34 ? stage1_inputData_0_delay_35_X : dataRam_0_io_rData_0_X);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_a_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_a_Y = (_zz_io_dataIn_0_payload_a_X_34 ? stage1_inputData_0_delay_35_Y : dataRam_0_io_rData_0_Y);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_a_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_a_Z = (_zz_io_dataIn_0_payload_a_X_34 ? stage1_inputData_0_delay_35_Z : dataRam_0_io_rData_0_Z);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_a_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_a_T = (_zz_io_dataIn_0_payload_a_X_34 ? stage1_inputData_0_delay_35_T : dataRam_0_io_rData_0_T);
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_b_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_b_X = pAddPort_0_s_delay_30_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_b_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_b_Y = pAddPort_0_s_delay_30_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_b_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_b_Z = pAddPort_0_s_delay_30_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_b_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_b_T = pAddPort_0_s_delay_30_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_0_payload_address = 17'bxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_0_payload_address = shiftRegs_addressOutFull_0_delay_30;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_valid = _zz_io_dataIn_1_valid_34;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_valid = _zz_io_dataIn_1_valid_64;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_valid = _zz_io_dataIn_1_valid_94;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_a_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_a_X = dataRam_0_io_rData_1_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_a_X = dataRam_0_io_rData_1_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_a_X = dataRam_0_io_rData_1_X;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_a_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_a_Y = dataRam_0_io_rData_1_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_a_Y = dataRam_0_io_rData_1_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_a_Y = dataRam_0_io_rData_1_Y;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_a_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_a_Z = dataRam_0_io_rData_1_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_a_Z = dataRam_0_io_rData_1_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_a_Z = dataRam_0_io_rData_1_Z;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_a_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_a_T = dataRam_0_io_rData_1_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_a_T = dataRam_0_io_rData_1_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_a_T = dataRam_0_io_rData_1_T;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_b_X = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_b_X = stage1_inputData_0_delay_35_X_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_b_X = pippenger_1_dataRam_0_io_rData_1_regNext_X;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_b_X = pippenger_1_dataRam_0_io_rData_1_regNext_X_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_b_Y = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_b_Y = stage1_inputData_0_delay_35_Y_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_b_Y = pippenger_1_dataRam_0_io_rData_1_regNext_Y;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_b_Y = pippenger_1_dataRam_0_io_rData_1_regNext_Y_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_b_Z = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_b_Z = stage1_inputData_0_delay_35_Z_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_b_Z = pippenger_1_dataRam_0_io_rData_1_regNext_Z;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_b_Z = pippenger_1_dataRam_0_io_rData_1_regNext_Z_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_b_T = 377'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_b_T = stage1_inputData_0_delay_35_T_1;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_b_T = pippenger_1_dataRam_0_io_rData_1_regNext_T;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_b_T = pippenger_1_dataRam_0_io_rData_1_regNext_T_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fifo_0_io_dataIn_1_payload_address = 17'bxxxxxxxxxxxxxxxxx;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        fifo_0_io_dataIn_1_payload_address = stage1_inputAddress_0_delay_35;
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        fifo_0_io_dataIn_1_payload_address = _zz_io_dataIn_1_payload_address_29;
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        fifo_0_io_dataIn_1_payload_address = {_zz_io_dataIn_1_payload_address_59,12'h001};
      end
      default : begin
      end
    endcase
  end

  assign io_dataOut_valid = outputValid;
  assign io_dataOut_payload_X = pAddPort_0_s_regNext_X;
  assign io_dataOut_payload_Y = pAddPort_0_s_regNext_Y;
  assign io_dataOut_payload_Z = pAddPort_0_s_regNext_Z;
  assign io_dataOut_payload_T = pAddPort_0_s_regNext_T;
  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    flushing_flushCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
        flushing_flushCnt_willIncrement = 1'b1;
      end
    endcase
  end

  assign flushing_flushCnt_willClear = 1'b0;
  assign flushing_flushCnt_willOverflow = (flushing_flushCnt_willOverflowIfInc && flushing_flushCnt_willIncrement);
  always @(*) begin
    if(flushing_flushCnt_willOverflow) begin
      flushing_flushCnt_valueNext = 17'h0;
    end else begin
      flushing_flushCnt_valueNext = (flushing_flushCnt_value + _zz_flushing_flushCnt_valueNext);
    end
    if(flushing_flushCnt_willClear) begin
      flushing_flushCnt_valueNext = 17'h0;
    end
  end

  always @(*) begin
    stage1_NCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          if(dataInBuffer_bufferOut_valid) begin
            if(stage1_GCnt_willOverflowIfInc) begin
              stage1_NCnt_willIncrement = 1'b1;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stage1_NCnt_willClear = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          if(dataInBuffer_bufferOut_valid) begin
            if(stage1_GCnt_willOverflowIfInc) begin
              if(dataInBuffer_bufferOut_payload_last) begin
                stage1_NCnt_willClear = 1'b1;
              end
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage1_NCnt_willOverflow = (stage1_NCnt_willOverflowIfInc && stage1_NCnt_willIncrement);
  always @(*) begin
    stage1_NCnt_valueNext = (stage1_NCnt_value + _zz_stage1_NCnt_valueNext);
    if(stage1_NCnt_willClear) begin
      stage1_NCnt_valueNext = 32'h0;
    end
  end

  always @(*) begin
    stage1_GCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(when_Pippenger_l153) begin
          if(dataInBuffer_bufferOut_valid) begin
            stage1_GCnt_willIncrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage1_GCnt_willClear = 1'b0;
  assign stage1_GCnt_willOverflow = (stage1_GCnt_willOverflowIfInc && stage1_GCnt_willIncrement);
  always @(*) begin
    if(stage1_GCnt_willOverflow) begin
      stage1_GCnt_valueNext = 5'h0;
    end else begin
      stage1_GCnt_valueNext = (stage1_GCnt_value + _zz_stage1_GCnt_valueNext);
    end
    if(stage1_GCnt_willClear) begin
      stage1_GCnt_valueNext = 5'h0;
    end
  end

  always @(*) begin
    stage1_emptyCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(!when_Pippenger_l153) begin
          if(!when_Pippenger_l168) begin
            stage1_emptyCnt_willIncrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    stage1_emptyCnt_willClear = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(!when_Pippenger_l153) begin
          if(when_Pippenger_l168) begin
            stage1_emptyCnt_willClear = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage1_emptyCnt_willOverflow = (stage1_emptyCnt_willOverflowIfInc && stage1_emptyCnt_willIncrement);
  always @(*) begin
    if(stage1_emptyCnt_willOverflow) begin
      stage1_emptyCnt_valueNext = 9'h0;
    end else begin
      stage1_emptyCnt_valueNext = (stage1_emptyCnt_value + _zz_stage1_emptyCnt_valueNext);
    end
    if(stage1_emptyCnt_willClear) begin
      stage1_emptyCnt_valueNext = 9'h0;
    end
  end

  assign stage1_inputBarrelID_0 = ({1'b0,_zz_stage1_inputBarrelID_0[12 : 0]} + _zz_stage1_inputBarrelID_0_1);
  assign _zz_stage1_inputBarrelIDAbs_0 = _zz__zz_stage1_inputBarrelIDAbs_0;
  assign stage1_inputBarrelIDAbs_0 = _zz_stage1_inputBarrelIDAbs_0_1[11:0];
  assign stage1_inputData_0_X = (_zz_stage1_inputData_0_X_5 ? pNegPort_n_X : dataInBuffer_bufferOut_payload_fragment_P_delay_6_X);
  assign stage1_inputData_0_Y = (_zz_stage1_inputData_0_X_5 ? pNegPort_n_Y : dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y);
  assign stage1_inputData_0_Z = (_zz_stage1_inputData_0_X_5 ? pNegPort_n_Z : dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z);
  assign stage1_inputData_0_T = (_zz_stage1_inputData_0_X_5 ? pNegPort_n_T : dataInBuffer_bufferOut_payload_fragment_P_delay_6_T);
  assign pAddPort_0_a_X = fifo_0_io_dataOut_payload_a_X;
  assign pAddPort_0_a_Y = fifo_0_io_dataOut_payload_a_Y;
  assign pAddPort_0_a_Z = fifo_0_io_dataOut_payload_a_Z;
  assign pAddPort_0_a_T = fifo_0_io_dataOut_payload_a_T;
  assign pAddPort_0_b_X = fifo_0_io_dataOut_payload_b_X;
  assign pAddPort_0_b_Y = fifo_0_io_dataOut_payload_b_Y;
  assign pAddPort_0_b_Z = fifo_0_io_dataOut_payload_b_Z;
  assign pAddPort_0_b_T = fifo_0_io_dataOut_payload_b_T;
  assign pNegPort_a_X = dataInBuffer_bufferOut_payload_fragment_P_X;
  assign pNegPort_a_Y = dataInBuffer_bufferOut_payload_fragment_P_Y;
  assign pNegPort_a_Z = dataInBuffer_bufferOut_payload_fragment_P_Z;
  assign pNegPort_a_T = dataInBuffer_bufferOut_payload_fragment_P_T;
  assign shiftRegs_validIn_0 = fifo_0_io_dataOut_valid;
  assign shiftRegs_addressIn_0 = fifo_0_io_dataOut_payload_address;
  always @(*) begin
    stage2_wCnt_willDecrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(!when_Pippenger_l207) begin
          if(stage2_waitCnt_willOverflowIfInc) begin
            stage2_wCnt_willDecrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage2_wCnt_willClear = 1'b0;
  assign stage2_wCnt_willUnderflow = (stage2_wCnt_willUnderflowIfDec && stage2_wCnt_willDecrement);
  always @(*) begin
    stage2_wCnt_valueNext = (stage2_wCnt_value - _zz_stage2_wCnt_valueNext);
    if(stage2_wCnt_willClear) begin
      stage2_wCnt_valueNext = 12'hfff;
    end
  end

  always @(*) begin
    stage2_GCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(when_Pippenger_l207) begin
          if(stage2_calCnt_willUnderflowIfDec) begin
            stage2_GCnt_willIncrement = 1'b1;
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage2_GCnt_willClear = 1'b0;
  assign stage2_GCnt_willOverflow = (stage2_GCnt_willOverflowIfInc && stage2_GCnt_willIncrement);
  always @(*) begin
    if(stage2_GCnt_willOverflow) begin
      stage2_GCnt_valueNext = 5'h0;
    end else begin
      stage2_GCnt_valueNext = (stage2_GCnt_value + _zz_stage2_GCnt_valueNext);
    end
    if(stage2_GCnt_willClear) begin
      stage2_GCnt_valueNext = 5'h0;
    end
  end

  always @(*) begin
    stage2_calCnt_willDecrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(when_Pippenger_l207) begin
          stage2_calCnt_willDecrement = 1'b1;
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage2_calCnt_willClear = 1'b0;
  assign stage2_calCnt_willUnderflow = (stage2_calCnt_willUnderflowIfDec && stage2_calCnt_willDecrement);
  always @(*) begin
    if(stage2_calCnt_willUnderflow) begin
      stage2_calCnt_valueNext = 2'b10;
    end else begin
      stage2_calCnt_valueNext = (stage2_calCnt_value - _zz_stage2_calCnt_valueNext);
    end
    if(stage2_calCnt_willClear) begin
      stage2_calCnt_valueNext = 2'b10;
    end
  end

  always @(*) begin
    stage2_waitCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(!when_Pippenger_l207) begin
          stage2_waitCnt_willIncrement = 1'b1;
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
      end
      default : begin
      end
    endcase
  end

  assign stage2_waitCnt_willClear = 1'b0;
  assign stage2_waitCnt_willOverflow = (stage2_waitCnt_willOverflowIfInc && stage2_waitCnt_willIncrement);
  always @(*) begin
    if(stage2_waitCnt_willOverflow) begin
      stage2_waitCnt_valueNext = 9'h0;
    end else begin
      stage2_waitCnt_valueNext = (stage2_waitCnt_value + _zz_stage2_waitCnt_valueNext);
    end
    if(stage2_waitCnt_willClear) begin
      stage2_waitCnt_valueNext = 9'h0;
    end
  end

  always @(*) begin
    stage3_GCnt_willDecrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(!when_Pippenger_l249) begin
          if(stage3_addWaitCnt_willOverflowIfInc) begin
            stage3_GCnt_willDecrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign stage3_GCnt_willClear = 1'b0;
  assign stage3_GCnt_willUnderflow = (stage3_GCnt_willUnderflowIfDec && stage3_GCnt_willDecrement);
  always @(*) begin
    if(stage3_GCnt_willUnderflow) begin
      stage3_GCnt_valueNext = 5'h13;
    end else begin
      stage3_GCnt_valueNext = (stage3_GCnt_value - _zz_stage3_GCnt_valueNext);
    end
    if(stage3_GCnt_willClear) begin
      stage3_GCnt_valueNext = 5'h13;
    end
  end

  always @(*) begin
    stage3_doubleCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(when_Pippenger_l249) begin
          if(stage3_doubleWaitCnt_willOverflowIfInc) begin
            stage3_doubleCnt_willIncrement = 1'b1;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign stage3_doubleCnt_willClear = 1'b0;
  assign stage3_doubleCnt_willOverflow = (stage3_doubleCnt_willOverflowIfInc && stage3_doubleCnt_willIncrement);
  always @(*) begin
    if(stage3_doubleCnt_willOverflow) begin
      stage3_doubleCnt_valueNext = 4'b0000;
    end else begin
      stage3_doubleCnt_valueNext = (stage3_doubleCnt_value + _zz_stage3_doubleCnt_valueNext);
    end
    if(stage3_doubleCnt_willClear) begin
      stage3_doubleCnt_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    stage3_doubleWaitCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(when_Pippenger_l249) begin
          stage3_doubleWaitCnt_willIncrement = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign stage3_doubleWaitCnt_willClear = 1'b0;
  assign stage3_doubleWaitCnt_willOverflow = (stage3_doubleWaitCnt_willOverflowIfInc && stage3_doubleWaitCnt_willIncrement);
  always @(*) begin
    if(stage3_doubleWaitCnt_willOverflow) begin
      stage3_doubleWaitCnt_valueNext = 9'h0;
    end else begin
      stage3_doubleWaitCnt_valueNext = (stage3_doubleWaitCnt_value + _zz_stage3_doubleWaitCnt_valueNext);
    end
    if(stage3_doubleWaitCnt_willClear) begin
      stage3_doubleWaitCnt_valueNext = 9'h0;
    end
  end

  always @(*) begin
    stage3_addWaitCnt_willIncrement = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(!when_Pippenger_l249) begin
          stage3_addWaitCnt_willIncrement = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign stage3_addWaitCnt_willClear = 1'b0;
  assign stage3_addWaitCnt_willOverflow = (stage3_addWaitCnt_willOverflowIfInc && stage3_addWaitCnt_willIncrement);
  always @(*) begin
    if(stage3_addWaitCnt_willOverflow) begin
      stage3_addWaitCnt_valueNext = 9'h0;
    end else begin
      stage3_addWaitCnt_valueNext = (stage3_addWaitCnt_value + _zz_stage3_addWaitCnt_valueNext);
    end
    if(stage3_addWaitCnt_willClear) begin
      stage3_addWaitCnt_valueNext = 9'h0;
    end
  end

  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
        if(!when_Pippenger_l153) begin
          if(!when_Pippenger_l168) begin
            if(stage1_emptyCnt_willOverflowIfInc) begin
              fsm_stateNext = fsm_enumDef_stage2;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
        if(!when_Pippenger_l207) begin
          if(stage2_waitCnt_willOverflowIfInc) begin
            if(stage2_wCnt_willUnderflowIfDec) begin
              fsm_stateNext = fsm_enumDef_stage3;
            end
          end
        end
      end
      (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
        if(!when_Pippenger_l249) begin
          if(stage3_addWaitCnt_willOverflowIfInc) begin
            if(stage3_GCnt_willUnderflowIfDec) begin
              fsm_stateNext = fsm_enumDef_stage1;
            end
          end
        end
      end
      default : begin
        if(flushing_flushCnt_willOverflowIfInc) begin
          fsm_stateNext = fsm_enumDef_stage1;
        end
      end
    endcase
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_flushing;
    end
  end

  assign when_Pippenger_l153 = (! stage1_waitReg);
  assign when_Pippenger_l168 = (fifo_0_io_dataOut_valid != 1'b0);
  assign when_Pippenger_l207 = (! stage2_waitReg);
  assign when_Pippenger_l249 = (! stage3_addReg);
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      dataInBuffer_validReg <= 1'b0;
      shiftRegs_validIn_delay_1_0 <= 1'b0;
      shiftRegs_validIn_delay_2_0 <= 1'b0;
      shiftRegs_validIn_delay_3_0 <= 1'b0;
      shiftRegs_validIn_delay_4_0 <= 1'b0;
      shiftRegs_validIn_delay_5_0 <= 1'b0;
      shiftRegs_validIn_delay_6_0 <= 1'b0;
      shiftRegs_validIn_delay_7_0 <= 1'b0;
      shiftRegs_validIn_delay_8_0 <= 1'b0;
      shiftRegs_validIn_delay_9_0 <= 1'b0;
      shiftRegs_validIn_delay_10_0 <= 1'b0;
      shiftRegs_validIn_delay_11_0 <= 1'b0;
      shiftRegs_validIn_delay_12_0 <= 1'b0;
      shiftRegs_validIn_delay_13_0 <= 1'b0;
      shiftRegs_validIn_delay_14_0 <= 1'b0;
      shiftRegs_validIn_delay_15_0 <= 1'b0;
      shiftRegs_validIn_delay_16_0 <= 1'b0;
      shiftRegs_validIn_delay_17_0 <= 1'b0;
      shiftRegs_validIn_delay_18_0 <= 1'b0;
      shiftRegs_validIn_delay_19_0 <= 1'b0;
      shiftRegs_validIn_delay_20_0 <= 1'b0;
      shiftRegs_validIn_delay_21_0 <= 1'b0;
      shiftRegs_validIn_delay_22_0 <= 1'b0;
      shiftRegs_validIn_delay_23_0 <= 1'b0;
      shiftRegs_validIn_delay_24_0 <= 1'b0;
      shiftRegs_validIn_delay_25_0 <= 1'b0;
      shiftRegs_validIn_delay_26_0 <= 1'b0;
      shiftRegs_validIn_delay_27_0 <= 1'b0;
      shiftRegs_validIn_delay_28_0 <= 1'b0;
      shiftRegs_validIn_delay_29_0 <= 1'b0;
      shiftRegs_validIn_delay_30_0 <= 1'b0;
      shiftRegs_validIn_delay_31_0 <= 1'b0;
      shiftRegs_validIn_delay_32_0 <= 1'b0;
      shiftRegs_validIn_delay_33_0 <= 1'b0;
      shiftRegs_validIn_delay_34_0 <= 1'b0;
      shiftRegs_validIn_delay_35_0 <= 1'b0;
      shiftRegs_validIn_delay_36_0 <= 1'b0;
      shiftRegs_validIn_delay_37_0 <= 1'b0;
      shiftRegs_validIn_delay_38_0 <= 1'b0;
      shiftRegs_validIn_delay_39_0 <= 1'b0;
      shiftRegs_validIn_delay_40_0 <= 1'b0;
      shiftRegs_validIn_delay_41_0 <= 1'b0;
      shiftRegs_validIn_delay_42_0 <= 1'b0;
      shiftRegs_validIn_delay_43_0 <= 1'b0;
      shiftRegs_validIn_delay_44_0 <= 1'b0;
      shiftRegs_validIn_delay_45_0 <= 1'b0;
      shiftRegs_validIn_delay_46_0 <= 1'b0;
      shiftRegs_validIn_delay_47_0 <= 1'b0;
      shiftRegs_validIn_delay_48_0 <= 1'b0;
      shiftRegs_validIn_delay_49_0 <= 1'b0;
      shiftRegs_validIn_delay_50_0 <= 1'b0;
      shiftRegs_validIn_delay_51_0 <= 1'b0;
      shiftRegs_validIn_delay_52_0 <= 1'b0;
      shiftRegs_validIn_delay_53_0 <= 1'b0;
      shiftRegs_validIn_delay_54_0 <= 1'b0;
      shiftRegs_validIn_delay_55_0 <= 1'b0;
      shiftRegs_validIn_delay_56_0 <= 1'b0;
      shiftRegs_validIn_delay_57_0 <= 1'b0;
      shiftRegs_validIn_delay_58_0 <= 1'b0;
      shiftRegs_validIn_delay_59_0 <= 1'b0;
      shiftRegs_validIn_delay_60_0 <= 1'b0;
      shiftRegs_validIn_delay_61_0 <= 1'b0;
      shiftRegs_validIn_delay_62_0 <= 1'b0;
      shiftRegs_validIn_delay_63_0 <= 1'b0;
      shiftRegs_validIn_delay_64_0 <= 1'b0;
      shiftRegs_validIn_delay_65_0 <= 1'b0;
      shiftRegs_validIn_delay_66_0 <= 1'b0;
      shiftRegs_validIn_delay_67_0 <= 1'b0;
      shiftRegs_validIn_delay_68_0 <= 1'b0;
      shiftRegs_validIn_delay_69_0 <= 1'b0;
      shiftRegs_validIn_delay_70_0 <= 1'b0;
      shiftRegs_validIn_delay_71_0 <= 1'b0;
      shiftRegs_validIn_delay_72_0 <= 1'b0;
      shiftRegs_validIn_delay_73_0 <= 1'b0;
      shiftRegs_validIn_delay_74_0 <= 1'b0;
      shiftRegs_validIn_delay_75_0 <= 1'b0;
      shiftRegs_validIn_delay_76_0 <= 1'b0;
      shiftRegs_validIn_delay_77_0 <= 1'b0;
      shiftRegs_validIn_delay_78_0 <= 1'b0;
      shiftRegs_validIn_delay_79_0 <= 1'b0;
      shiftRegs_validIn_delay_80_0 <= 1'b0;
      shiftRegs_validIn_delay_81_0 <= 1'b0;
      shiftRegs_validIn_delay_82_0 <= 1'b0;
      shiftRegs_validIn_delay_83_0 <= 1'b0;
      shiftRegs_validIn_delay_84_0 <= 1'b0;
      shiftRegs_validIn_delay_85_0 <= 1'b0;
      shiftRegs_validIn_delay_86_0 <= 1'b0;
      shiftRegs_validIn_delay_87_0 <= 1'b0;
      shiftRegs_validIn_delay_88_0 <= 1'b0;
      shiftRegs_validIn_delay_89_0 <= 1'b0;
      shiftRegs_validIn_delay_90_0 <= 1'b0;
      shiftRegs_validIn_delay_91_0 <= 1'b0;
      shiftRegs_validIn_delay_92_0 <= 1'b0;
      shiftRegs_validIn_delay_93_0 <= 1'b0;
      shiftRegs_validIn_delay_94_0 <= 1'b0;
      shiftRegs_validIn_delay_95_0 <= 1'b0;
      shiftRegs_validIn_delay_96_0 <= 1'b0;
      shiftRegs_validIn_delay_97_0 <= 1'b0;
      shiftRegs_validIn_delay_98_0 <= 1'b0;
      shiftRegs_validIn_delay_99_0 <= 1'b0;
      shiftRegs_validIn_delay_100_0 <= 1'b0;
      shiftRegs_validIn_delay_101_0 <= 1'b0;
      shiftRegs_validIn_delay_102_0 <= 1'b0;
      shiftRegs_validIn_delay_103_0 <= 1'b0;
      shiftRegs_validIn_delay_104_0 <= 1'b0;
      shiftRegs_validIn_delay_105_0 <= 1'b0;
      shiftRegs_validIn_delay_106_0 <= 1'b0;
      shiftRegs_validIn_delay_107_0 <= 1'b0;
      shiftRegs_validIn_delay_108_0 <= 1'b0;
      shiftRegs_validIn_delay_109_0 <= 1'b0;
      shiftRegs_validIn_delay_110_0 <= 1'b0;
      shiftRegs_validIn_delay_111_0 <= 1'b0;
      shiftRegs_validIn_delay_112_0 <= 1'b0;
      shiftRegs_validIn_delay_113_0 <= 1'b0;
      shiftRegs_validIn_delay_114_0 <= 1'b0;
      shiftRegs_validIn_delay_115_0 <= 1'b0;
      shiftRegs_validIn_delay_116_0 <= 1'b0;
      shiftRegs_validIn_delay_117_0 <= 1'b0;
      shiftRegs_validIn_delay_118_0 <= 1'b0;
      shiftRegs_validIn_delay_119_0 <= 1'b0;
      shiftRegs_validIn_delay_120_0 <= 1'b0;
      shiftRegs_validIn_delay_121_0 <= 1'b0;
      shiftRegs_validIn_delay_122_0 <= 1'b0;
      shiftRegs_validIn_delay_123_0 <= 1'b0;
      shiftRegs_validIn_delay_124_0 <= 1'b0;
      shiftRegs_validIn_delay_125_0 <= 1'b0;
      shiftRegs_validIn_delay_126_0 <= 1'b0;
      shiftRegs_validIn_delay_127_0 <= 1'b0;
      shiftRegs_validIn_delay_128_0 <= 1'b0;
      shiftRegs_validIn_delay_129_0 <= 1'b0;
      shiftRegs_validIn_delay_130_0 <= 1'b0;
      shiftRegs_validIn_delay_131_0 <= 1'b0;
      shiftRegs_validIn_delay_132_0 <= 1'b0;
      shiftRegs_validIn_delay_133_0 <= 1'b0;
      shiftRegs_validIn_delay_134_0 <= 1'b0;
      shiftRegs_validIn_delay_135_0 <= 1'b0;
      shiftRegs_validIn_delay_136_0 <= 1'b0;
      shiftRegs_validIn_delay_137_0 <= 1'b0;
      shiftRegs_validIn_delay_138_0 <= 1'b0;
      shiftRegs_validIn_delay_139_0 <= 1'b0;
      shiftRegs_validIn_delay_140_0 <= 1'b0;
      shiftRegs_validIn_delay_141_0 <= 1'b0;
      shiftRegs_validIn_delay_142_0 <= 1'b0;
      shiftRegs_validIn_delay_143_0 <= 1'b0;
      shiftRegs_validIn_delay_144_0 <= 1'b0;
      shiftRegs_validIn_delay_145_0 <= 1'b0;
      shiftRegs_validIn_delay_146_0 <= 1'b0;
      shiftRegs_validIn_delay_147_0 <= 1'b0;
      shiftRegs_validIn_delay_148_0 <= 1'b0;
      shiftRegs_validIn_delay_149_0 <= 1'b0;
      shiftRegs_validIn_delay_150_0 <= 1'b0;
      shiftRegs_validIn_delay_151_0 <= 1'b0;
      shiftRegs_validIn_delay_152_0 <= 1'b0;
      shiftRegs_validIn_delay_153_0 <= 1'b0;
      shiftRegs_validIn_delay_154_0 <= 1'b0;
      shiftRegs_validIn_delay_155_0 <= 1'b0;
      shiftRegs_validIn_delay_156_0 <= 1'b0;
      shiftRegs_validIn_delay_157_0 <= 1'b0;
      shiftRegs_validIn_delay_158_0 <= 1'b0;
      shiftRegs_validIn_delay_159_0 <= 1'b0;
      shiftRegs_validIn_delay_160_0 <= 1'b0;
      shiftRegs_validIn_delay_161_0 <= 1'b0;
      shiftRegs_validIn_delay_162_0 <= 1'b0;
      shiftRegs_validIn_delay_163_0 <= 1'b0;
      shiftRegs_validIn_delay_164_0 <= 1'b0;
      shiftRegs_validIn_delay_165_0 <= 1'b0;
      shiftRegs_validIn_delay_166_0 <= 1'b0;
      shiftRegs_validIn_delay_167_0 <= 1'b0;
      shiftRegs_validIn_delay_168_0 <= 1'b0;
      shiftRegs_validIn_delay_169_0 <= 1'b0;
      shiftRegs_validIn_delay_170_0 <= 1'b0;
      shiftRegs_validIn_delay_171_0 <= 1'b0;
      shiftRegs_validIn_delay_172_0 <= 1'b0;
      shiftRegs_validIn_delay_173_0 <= 1'b0;
      shiftRegs_validIn_delay_174_0 <= 1'b0;
      shiftRegs_validIn_delay_175_0 <= 1'b0;
      shiftRegs_validIn_delay_176_0 <= 1'b0;
      shiftRegs_validIn_delay_177_0 <= 1'b0;
      shiftRegs_validIn_delay_178_0 <= 1'b0;
      shiftRegs_validIn_delay_179_0 <= 1'b0;
      shiftRegs_validIn_delay_180_0 <= 1'b0;
      shiftRegs_validIn_delay_181_0 <= 1'b0;
      shiftRegs_validIn_delay_182_0 <= 1'b0;
      shiftRegs_validIn_delay_183_0 <= 1'b0;
      shiftRegs_validIn_delay_184_0 <= 1'b0;
      shiftRegs_validIn_delay_185_0 <= 1'b0;
      shiftRegs_validIn_delay_186_0 <= 1'b0;
      shiftRegs_validIn_delay_187_0 <= 1'b0;
      shiftRegs_validIn_delay_188_0 <= 1'b0;
      shiftRegs_validIn_delay_189_0 <= 1'b0;
      shiftRegs_validIn_delay_190_0 <= 1'b0;
      shiftRegs_validIn_delay_191_0 <= 1'b0;
      shiftRegs_validIn_delay_192_0 <= 1'b0;
      shiftRegs_validIn_delay_193_0 <= 1'b0;
      shiftRegs_validIn_delay_194_0 <= 1'b0;
      shiftRegs_validIn_delay_195_0 <= 1'b0;
      shiftRegs_validIn_delay_196_0 <= 1'b0;
      shiftRegs_validIn_delay_197_0 <= 1'b0;
      shiftRegs_validIn_delay_198_0 <= 1'b0;
      shiftRegs_validIn_delay_199_0 <= 1'b0;
      shiftRegs_validIn_delay_200_0 <= 1'b0;
      shiftRegs_validIn_delay_201_0 <= 1'b0;
      shiftRegs_validIn_delay_202_0 <= 1'b0;
      shiftRegs_validIn_delay_203_0 <= 1'b0;
      shiftRegs_validIn_delay_204_0 <= 1'b0;
      shiftRegs_validIn_delay_205_0 <= 1'b0;
      shiftRegs_validIn_delay_206_0 <= 1'b0;
      shiftRegs_validIn_delay_207_0 <= 1'b0;
      shiftRegs_validIn_delay_208_0 <= 1'b0;
      shiftRegs_validIn_delay_209_0 <= 1'b0;
      shiftRegs_validIn_delay_210_0 <= 1'b0;
      shiftRegs_validIn_delay_211_0 <= 1'b0;
      shiftRegs_validIn_delay_212_0 <= 1'b0;
      shiftRegs_validIn_delay_213_0 <= 1'b0;
      shiftRegs_validIn_delay_214_0 <= 1'b0;
      shiftRegs_validIn_delay_215_0 <= 1'b0;
      shiftRegs_validIn_delay_216_0 <= 1'b0;
      shiftRegs_validIn_delay_217_0 <= 1'b0;
      shiftRegs_validIn_delay_218_0 <= 1'b0;
      shiftRegs_validIn_delay_219_0 <= 1'b0;
      shiftRegs_validIn_delay_220_0 <= 1'b0;
      shiftRegs_validIn_delay_221_0 <= 1'b0;
      shiftRegs_validIn_delay_222_0 <= 1'b0;
      shiftRegs_validIn_delay_223_0 <= 1'b0;
      shiftRegs_validIn_delay_224_0 <= 1'b0;
      shiftRegs_validIn_delay_225_0 <= 1'b0;
      shiftRegs_validIn_delay_226_0 <= 1'b0;
      shiftRegs_validIn_delay_227_0 <= 1'b0;
      shiftRegs_validIn_delay_228_0 <= 1'b0;
      shiftRegs_validIn_delay_229_0 <= 1'b0;
      shiftRegs_validIn_delay_230_0 <= 1'b0;
      shiftRegs_validIn_delay_231_0 <= 1'b0;
      shiftRegs_validIn_delay_232_0 <= 1'b0;
      shiftRegs_validIn_delay_233_0 <= 1'b0;
      shiftRegs_validIn_delay_234_0 <= 1'b0;
      shiftRegs_validIn_delay_235_0 <= 1'b0;
      shiftRegs_validIn_delay_236_0 <= 1'b0;
      shiftRegs_validIn_delay_237_0 <= 1'b0;
      shiftRegs_validIn_delay_238_0 <= 1'b0;
      shiftRegs_validIn_delay_239_0 <= 1'b0;
      shiftRegs_validIn_delay_240_0 <= 1'b0;
      shiftRegs_validIn_delay_241_0 <= 1'b0;
      shiftRegs_validIn_delay_242_0 <= 1'b0;
      shiftRegs_validIn_delay_243_0 <= 1'b0;
      shiftRegs_validIn_delay_244_0 <= 1'b0;
      shiftRegs_validIn_delay_245_0 <= 1'b0;
      shiftRegs_validIn_delay_246_0 <= 1'b0;
      shiftRegs_validIn_delay_247_0 <= 1'b0;
      shiftRegs_validIn_delay_248_0 <= 1'b0;
      shiftRegs_validIn_delay_249_0 <= 1'b0;
      shiftRegs_validIn_delay_250_0 <= 1'b0;
      shiftRegs_validIn_delay_251_0 <= 1'b0;
      shiftRegs_validIn_delay_252_0 <= 1'b0;
      shiftRegs_validIn_delay_253_0 <= 1'b0;
      shiftRegs_validIn_delay_254_0 <= 1'b0;
      shiftRegs_validOut_0 <= 1'b0;
      shiftRegs_validOut_delay_1_0 <= 1'b0;
      shiftRegs_validOut_delay_2_0 <= 1'b0;
      shiftRegs_validOut_delay_3_0 <= 1'b0;
      shiftRegs_validOut_delay_4_0 <= 1'b0;
      shiftRegs_validOutFull_0 <= 1'b0;
      outputValid <= 1'b0;
      flushing_flushCnt_value <= 17'h0;
      flushing_flushCnt_willOverflowIfInc <= 1'b0;
      stage1_NCnt_value <= 32'h0;
      stage1_NCnt_willOverflowIfInc <= 1'b0;
      stage1_GCnt_value <= 5'h0;
      stage1_GCnt_willOverflowIfInc <= 1'b0;
      stage1_waitReg <= 1'b0;
      stage1_emptyCnt_value <= 9'h0;
      stage1_emptyCnt_willOverflowIfInc <= 1'b0;
      stage1_needAdd1_0 <= 1'b0;
      _zz_stage1_inputValid_0 <= 1'b0;
      _zz_stage1_inputValid_0_1 <= 1'b0;
      _zz_stage1_inputValid_0_2 <= 1'b0;
      _zz_stage1_inputValid_0_3 <= 1'b0;
      _zz_stage1_inputValid_0_4 <= 1'b0;
      stage1_inputValid_0 <= 1'b0;
      stage2_wCnt_value <= 12'hfff;
      stage2_wCnt_willUnderflowIfDec <= 1'b0;
      stage2_GCnt_value <= 5'h0;
      stage2_GCnt_willOverflowIfInc <= 1'b0;
      stage2_calCnt_value <= 2'b10;
      stage2_calCnt_willUnderflowIfDec <= 1'b0;
      stage2_waitReg <= 1'b0;
      stage2_waitCnt_value <= 9'h0;
      stage2_waitCnt_willOverflowIfInc <= 1'b0;
      stage3_GCnt_value <= 5'h13;
      stage3_GCnt_willUnderflowIfDec <= 1'b0;
      stage3_doubleCnt_value <= 4'b0000;
      stage3_doubleCnt_willOverflowIfInc <= 1'b0;
      stage3_doubleWaitCnt_value <= 9'h0;
      stage3_doubleWaitCnt_willOverflowIfInc <= 1'b0;
      stage3_addReg <= 1'b0;
      stage3_addWaitCnt_value <= 9'h0;
      stage3_addWaitCnt_willOverflowIfInc <= 1'b0;
      fsm_stateReg <= fsm_enumDef_flushing;
    end else begin
      if(io_dataIn_valid) begin
        dataInBuffer_validReg <= 1'b1;
      end else begin
        if(dataInBuffer_bufferOut_ready) begin
          dataInBuffer_validReg <= 1'b0;
        end
      end
      shiftRegs_validIn_delay_1_0 <= shiftRegs_validIn_0;
      shiftRegs_validIn_delay_2_0 <= shiftRegs_validIn_delay_1_0;
      shiftRegs_validIn_delay_3_0 <= shiftRegs_validIn_delay_2_0;
      shiftRegs_validIn_delay_4_0 <= shiftRegs_validIn_delay_3_0;
      shiftRegs_validIn_delay_5_0 <= shiftRegs_validIn_delay_4_0;
      shiftRegs_validIn_delay_6_0 <= shiftRegs_validIn_delay_5_0;
      shiftRegs_validIn_delay_7_0 <= shiftRegs_validIn_delay_6_0;
      shiftRegs_validIn_delay_8_0 <= shiftRegs_validIn_delay_7_0;
      shiftRegs_validIn_delay_9_0 <= shiftRegs_validIn_delay_8_0;
      shiftRegs_validIn_delay_10_0 <= shiftRegs_validIn_delay_9_0;
      shiftRegs_validIn_delay_11_0 <= shiftRegs_validIn_delay_10_0;
      shiftRegs_validIn_delay_12_0 <= shiftRegs_validIn_delay_11_0;
      shiftRegs_validIn_delay_13_0 <= shiftRegs_validIn_delay_12_0;
      shiftRegs_validIn_delay_14_0 <= shiftRegs_validIn_delay_13_0;
      shiftRegs_validIn_delay_15_0 <= shiftRegs_validIn_delay_14_0;
      shiftRegs_validIn_delay_16_0 <= shiftRegs_validIn_delay_15_0;
      shiftRegs_validIn_delay_17_0 <= shiftRegs_validIn_delay_16_0;
      shiftRegs_validIn_delay_18_0 <= shiftRegs_validIn_delay_17_0;
      shiftRegs_validIn_delay_19_0 <= shiftRegs_validIn_delay_18_0;
      shiftRegs_validIn_delay_20_0 <= shiftRegs_validIn_delay_19_0;
      shiftRegs_validIn_delay_21_0 <= shiftRegs_validIn_delay_20_0;
      shiftRegs_validIn_delay_22_0 <= shiftRegs_validIn_delay_21_0;
      shiftRegs_validIn_delay_23_0 <= shiftRegs_validIn_delay_22_0;
      shiftRegs_validIn_delay_24_0 <= shiftRegs_validIn_delay_23_0;
      shiftRegs_validIn_delay_25_0 <= shiftRegs_validIn_delay_24_0;
      shiftRegs_validIn_delay_26_0 <= shiftRegs_validIn_delay_25_0;
      shiftRegs_validIn_delay_27_0 <= shiftRegs_validIn_delay_26_0;
      shiftRegs_validIn_delay_28_0 <= shiftRegs_validIn_delay_27_0;
      shiftRegs_validIn_delay_29_0 <= shiftRegs_validIn_delay_28_0;
      shiftRegs_validIn_delay_30_0 <= shiftRegs_validIn_delay_29_0;
      shiftRegs_validIn_delay_31_0 <= shiftRegs_validIn_delay_30_0;
      shiftRegs_validIn_delay_32_0 <= shiftRegs_validIn_delay_31_0;
      shiftRegs_validIn_delay_33_0 <= shiftRegs_validIn_delay_32_0;
      shiftRegs_validIn_delay_34_0 <= shiftRegs_validIn_delay_33_0;
      shiftRegs_validIn_delay_35_0 <= shiftRegs_validIn_delay_34_0;
      shiftRegs_validIn_delay_36_0 <= shiftRegs_validIn_delay_35_0;
      shiftRegs_validIn_delay_37_0 <= shiftRegs_validIn_delay_36_0;
      shiftRegs_validIn_delay_38_0 <= shiftRegs_validIn_delay_37_0;
      shiftRegs_validIn_delay_39_0 <= shiftRegs_validIn_delay_38_0;
      shiftRegs_validIn_delay_40_0 <= shiftRegs_validIn_delay_39_0;
      shiftRegs_validIn_delay_41_0 <= shiftRegs_validIn_delay_40_0;
      shiftRegs_validIn_delay_42_0 <= shiftRegs_validIn_delay_41_0;
      shiftRegs_validIn_delay_43_0 <= shiftRegs_validIn_delay_42_0;
      shiftRegs_validIn_delay_44_0 <= shiftRegs_validIn_delay_43_0;
      shiftRegs_validIn_delay_45_0 <= shiftRegs_validIn_delay_44_0;
      shiftRegs_validIn_delay_46_0 <= shiftRegs_validIn_delay_45_0;
      shiftRegs_validIn_delay_47_0 <= shiftRegs_validIn_delay_46_0;
      shiftRegs_validIn_delay_48_0 <= shiftRegs_validIn_delay_47_0;
      shiftRegs_validIn_delay_49_0 <= shiftRegs_validIn_delay_48_0;
      shiftRegs_validIn_delay_50_0 <= shiftRegs_validIn_delay_49_0;
      shiftRegs_validIn_delay_51_0 <= shiftRegs_validIn_delay_50_0;
      shiftRegs_validIn_delay_52_0 <= shiftRegs_validIn_delay_51_0;
      shiftRegs_validIn_delay_53_0 <= shiftRegs_validIn_delay_52_0;
      shiftRegs_validIn_delay_54_0 <= shiftRegs_validIn_delay_53_0;
      shiftRegs_validIn_delay_55_0 <= shiftRegs_validIn_delay_54_0;
      shiftRegs_validIn_delay_56_0 <= shiftRegs_validIn_delay_55_0;
      shiftRegs_validIn_delay_57_0 <= shiftRegs_validIn_delay_56_0;
      shiftRegs_validIn_delay_58_0 <= shiftRegs_validIn_delay_57_0;
      shiftRegs_validIn_delay_59_0 <= shiftRegs_validIn_delay_58_0;
      shiftRegs_validIn_delay_60_0 <= shiftRegs_validIn_delay_59_0;
      shiftRegs_validIn_delay_61_0 <= shiftRegs_validIn_delay_60_0;
      shiftRegs_validIn_delay_62_0 <= shiftRegs_validIn_delay_61_0;
      shiftRegs_validIn_delay_63_0 <= shiftRegs_validIn_delay_62_0;
      shiftRegs_validIn_delay_64_0 <= shiftRegs_validIn_delay_63_0;
      shiftRegs_validIn_delay_65_0 <= shiftRegs_validIn_delay_64_0;
      shiftRegs_validIn_delay_66_0 <= shiftRegs_validIn_delay_65_0;
      shiftRegs_validIn_delay_67_0 <= shiftRegs_validIn_delay_66_0;
      shiftRegs_validIn_delay_68_0 <= shiftRegs_validIn_delay_67_0;
      shiftRegs_validIn_delay_69_0 <= shiftRegs_validIn_delay_68_0;
      shiftRegs_validIn_delay_70_0 <= shiftRegs_validIn_delay_69_0;
      shiftRegs_validIn_delay_71_0 <= shiftRegs_validIn_delay_70_0;
      shiftRegs_validIn_delay_72_0 <= shiftRegs_validIn_delay_71_0;
      shiftRegs_validIn_delay_73_0 <= shiftRegs_validIn_delay_72_0;
      shiftRegs_validIn_delay_74_0 <= shiftRegs_validIn_delay_73_0;
      shiftRegs_validIn_delay_75_0 <= shiftRegs_validIn_delay_74_0;
      shiftRegs_validIn_delay_76_0 <= shiftRegs_validIn_delay_75_0;
      shiftRegs_validIn_delay_77_0 <= shiftRegs_validIn_delay_76_0;
      shiftRegs_validIn_delay_78_0 <= shiftRegs_validIn_delay_77_0;
      shiftRegs_validIn_delay_79_0 <= shiftRegs_validIn_delay_78_0;
      shiftRegs_validIn_delay_80_0 <= shiftRegs_validIn_delay_79_0;
      shiftRegs_validIn_delay_81_0 <= shiftRegs_validIn_delay_80_0;
      shiftRegs_validIn_delay_82_0 <= shiftRegs_validIn_delay_81_0;
      shiftRegs_validIn_delay_83_0 <= shiftRegs_validIn_delay_82_0;
      shiftRegs_validIn_delay_84_0 <= shiftRegs_validIn_delay_83_0;
      shiftRegs_validIn_delay_85_0 <= shiftRegs_validIn_delay_84_0;
      shiftRegs_validIn_delay_86_0 <= shiftRegs_validIn_delay_85_0;
      shiftRegs_validIn_delay_87_0 <= shiftRegs_validIn_delay_86_0;
      shiftRegs_validIn_delay_88_0 <= shiftRegs_validIn_delay_87_0;
      shiftRegs_validIn_delay_89_0 <= shiftRegs_validIn_delay_88_0;
      shiftRegs_validIn_delay_90_0 <= shiftRegs_validIn_delay_89_0;
      shiftRegs_validIn_delay_91_0 <= shiftRegs_validIn_delay_90_0;
      shiftRegs_validIn_delay_92_0 <= shiftRegs_validIn_delay_91_0;
      shiftRegs_validIn_delay_93_0 <= shiftRegs_validIn_delay_92_0;
      shiftRegs_validIn_delay_94_0 <= shiftRegs_validIn_delay_93_0;
      shiftRegs_validIn_delay_95_0 <= shiftRegs_validIn_delay_94_0;
      shiftRegs_validIn_delay_96_0 <= shiftRegs_validIn_delay_95_0;
      shiftRegs_validIn_delay_97_0 <= shiftRegs_validIn_delay_96_0;
      shiftRegs_validIn_delay_98_0 <= shiftRegs_validIn_delay_97_0;
      shiftRegs_validIn_delay_99_0 <= shiftRegs_validIn_delay_98_0;
      shiftRegs_validIn_delay_100_0 <= shiftRegs_validIn_delay_99_0;
      shiftRegs_validIn_delay_101_0 <= shiftRegs_validIn_delay_100_0;
      shiftRegs_validIn_delay_102_0 <= shiftRegs_validIn_delay_101_0;
      shiftRegs_validIn_delay_103_0 <= shiftRegs_validIn_delay_102_0;
      shiftRegs_validIn_delay_104_0 <= shiftRegs_validIn_delay_103_0;
      shiftRegs_validIn_delay_105_0 <= shiftRegs_validIn_delay_104_0;
      shiftRegs_validIn_delay_106_0 <= shiftRegs_validIn_delay_105_0;
      shiftRegs_validIn_delay_107_0 <= shiftRegs_validIn_delay_106_0;
      shiftRegs_validIn_delay_108_0 <= shiftRegs_validIn_delay_107_0;
      shiftRegs_validIn_delay_109_0 <= shiftRegs_validIn_delay_108_0;
      shiftRegs_validIn_delay_110_0 <= shiftRegs_validIn_delay_109_0;
      shiftRegs_validIn_delay_111_0 <= shiftRegs_validIn_delay_110_0;
      shiftRegs_validIn_delay_112_0 <= shiftRegs_validIn_delay_111_0;
      shiftRegs_validIn_delay_113_0 <= shiftRegs_validIn_delay_112_0;
      shiftRegs_validIn_delay_114_0 <= shiftRegs_validIn_delay_113_0;
      shiftRegs_validIn_delay_115_0 <= shiftRegs_validIn_delay_114_0;
      shiftRegs_validIn_delay_116_0 <= shiftRegs_validIn_delay_115_0;
      shiftRegs_validIn_delay_117_0 <= shiftRegs_validIn_delay_116_0;
      shiftRegs_validIn_delay_118_0 <= shiftRegs_validIn_delay_117_0;
      shiftRegs_validIn_delay_119_0 <= shiftRegs_validIn_delay_118_0;
      shiftRegs_validIn_delay_120_0 <= shiftRegs_validIn_delay_119_0;
      shiftRegs_validIn_delay_121_0 <= shiftRegs_validIn_delay_120_0;
      shiftRegs_validIn_delay_122_0 <= shiftRegs_validIn_delay_121_0;
      shiftRegs_validIn_delay_123_0 <= shiftRegs_validIn_delay_122_0;
      shiftRegs_validIn_delay_124_0 <= shiftRegs_validIn_delay_123_0;
      shiftRegs_validIn_delay_125_0 <= shiftRegs_validIn_delay_124_0;
      shiftRegs_validIn_delay_126_0 <= shiftRegs_validIn_delay_125_0;
      shiftRegs_validIn_delay_127_0 <= shiftRegs_validIn_delay_126_0;
      shiftRegs_validIn_delay_128_0 <= shiftRegs_validIn_delay_127_0;
      shiftRegs_validIn_delay_129_0 <= shiftRegs_validIn_delay_128_0;
      shiftRegs_validIn_delay_130_0 <= shiftRegs_validIn_delay_129_0;
      shiftRegs_validIn_delay_131_0 <= shiftRegs_validIn_delay_130_0;
      shiftRegs_validIn_delay_132_0 <= shiftRegs_validIn_delay_131_0;
      shiftRegs_validIn_delay_133_0 <= shiftRegs_validIn_delay_132_0;
      shiftRegs_validIn_delay_134_0 <= shiftRegs_validIn_delay_133_0;
      shiftRegs_validIn_delay_135_0 <= shiftRegs_validIn_delay_134_0;
      shiftRegs_validIn_delay_136_0 <= shiftRegs_validIn_delay_135_0;
      shiftRegs_validIn_delay_137_0 <= shiftRegs_validIn_delay_136_0;
      shiftRegs_validIn_delay_138_0 <= shiftRegs_validIn_delay_137_0;
      shiftRegs_validIn_delay_139_0 <= shiftRegs_validIn_delay_138_0;
      shiftRegs_validIn_delay_140_0 <= shiftRegs_validIn_delay_139_0;
      shiftRegs_validIn_delay_141_0 <= shiftRegs_validIn_delay_140_0;
      shiftRegs_validIn_delay_142_0 <= shiftRegs_validIn_delay_141_0;
      shiftRegs_validIn_delay_143_0 <= shiftRegs_validIn_delay_142_0;
      shiftRegs_validIn_delay_144_0 <= shiftRegs_validIn_delay_143_0;
      shiftRegs_validIn_delay_145_0 <= shiftRegs_validIn_delay_144_0;
      shiftRegs_validIn_delay_146_0 <= shiftRegs_validIn_delay_145_0;
      shiftRegs_validIn_delay_147_0 <= shiftRegs_validIn_delay_146_0;
      shiftRegs_validIn_delay_148_0 <= shiftRegs_validIn_delay_147_0;
      shiftRegs_validIn_delay_149_0 <= shiftRegs_validIn_delay_148_0;
      shiftRegs_validIn_delay_150_0 <= shiftRegs_validIn_delay_149_0;
      shiftRegs_validIn_delay_151_0 <= shiftRegs_validIn_delay_150_0;
      shiftRegs_validIn_delay_152_0 <= shiftRegs_validIn_delay_151_0;
      shiftRegs_validIn_delay_153_0 <= shiftRegs_validIn_delay_152_0;
      shiftRegs_validIn_delay_154_0 <= shiftRegs_validIn_delay_153_0;
      shiftRegs_validIn_delay_155_0 <= shiftRegs_validIn_delay_154_0;
      shiftRegs_validIn_delay_156_0 <= shiftRegs_validIn_delay_155_0;
      shiftRegs_validIn_delay_157_0 <= shiftRegs_validIn_delay_156_0;
      shiftRegs_validIn_delay_158_0 <= shiftRegs_validIn_delay_157_0;
      shiftRegs_validIn_delay_159_0 <= shiftRegs_validIn_delay_158_0;
      shiftRegs_validIn_delay_160_0 <= shiftRegs_validIn_delay_159_0;
      shiftRegs_validIn_delay_161_0 <= shiftRegs_validIn_delay_160_0;
      shiftRegs_validIn_delay_162_0 <= shiftRegs_validIn_delay_161_0;
      shiftRegs_validIn_delay_163_0 <= shiftRegs_validIn_delay_162_0;
      shiftRegs_validIn_delay_164_0 <= shiftRegs_validIn_delay_163_0;
      shiftRegs_validIn_delay_165_0 <= shiftRegs_validIn_delay_164_0;
      shiftRegs_validIn_delay_166_0 <= shiftRegs_validIn_delay_165_0;
      shiftRegs_validIn_delay_167_0 <= shiftRegs_validIn_delay_166_0;
      shiftRegs_validIn_delay_168_0 <= shiftRegs_validIn_delay_167_0;
      shiftRegs_validIn_delay_169_0 <= shiftRegs_validIn_delay_168_0;
      shiftRegs_validIn_delay_170_0 <= shiftRegs_validIn_delay_169_0;
      shiftRegs_validIn_delay_171_0 <= shiftRegs_validIn_delay_170_0;
      shiftRegs_validIn_delay_172_0 <= shiftRegs_validIn_delay_171_0;
      shiftRegs_validIn_delay_173_0 <= shiftRegs_validIn_delay_172_0;
      shiftRegs_validIn_delay_174_0 <= shiftRegs_validIn_delay_173_0;
      shiftRegs_validIn_delay_175_0 <= shiftRegs_validIn_delay_174_0;
      shiftRegs_validIn_delay_176_0 <= shiftRegs_validIn_delay_175_0;
      shiftRegs_validIn_delay_177_0 <= shiftRegs_validIn_delay_176_0;
      shiftRegs_validIn_delay_178_0 <= shiftRegs_validIn_delay_177_0;
      shiftRegs_validIn_delay_179_0 <= shiftRegs_validIn_delay_178_0;
      shiftRegs_validIn_delay_180_0 <= shiftRegs_validIn_delay_179_0;
      shiftRegs_validIn_delay_181_0 <= shiftRegs_validIn_delay_180_0;
      shiftRegs_validIn_delay_182_0 <= shiftRegs_validIn_delay_181_0;
      shiftRegs_validIn_delay_183_0 <= shiftRegs_validIn_delay_182_0;
      shiftRegs_validIn_delay_184_0 <= shiftRegs_validIn_delay_183_0;
      shiftRegs_validIn_delay_185_0 <= shiftRegs_validIn_delay_184_0;
      shiftRegs_validIn_delay_186_0 <= shiftRegs_validIn_delay_185_0;
      shiftRegs_validIn_delay_187_0 <= shiftRegs_validIn_delay_186_0;
      shiftRegs_validIn_delay_188_0 <= shiftRegs_validIn_delay_187_0;
      shiftRegs_validIn_delay_189_0 <= shiftRegs_validIn_delay_188_0;
      shiftRegs_validIn_delay_190_0 <= shiftRegs_validIn_delay_189_0;
      shiftRegs_validIn_delay_191_0 <= shiftRegs_validIn_delay_190_0;
      shiftRegs_validIn_delay_192_0 <= shiftRegs_validIn_delay_191_0;
      shiftRegs_validIn_delay_193_0 <= shiftRegs_validIn_delay_192_0;
      shiftRegs_validIn_delay_194_0 <= shiftRegs_validIn_delay_193_0;
      shiftRegs_validIn_delay_195_0 <= shiftRegs_validIn_delay_194_0;
      shiftRegs_validIn_delay_196_0 <= shiftRegs_validIn_delay_195_0;
      shiftRegs_validIn_delay_197_0 <= shiftRegs_validIn_delay_196_0;
      shiftRegs_validIn_delay_198_0 <= shiftRegs_validIn_delay_197_0;
      shiftRegs_validIn_delay_199_0 <= shiftRegs_validIn_delay_198_0;
      shiftRegs_validIn_delay_200_0 <= shiftRegs_validIn_delay_199_0;
      shiftRegs_validIn_delay_201_0 <= shiftRegs_validIn_delay_200_0;
      shiftRegs_validIn_delay_202_0 <= shiftRegs_validIn_delay_201_0;
      shiftRegs_validIn_delay_203_0 <= shiftRegs_validIn_delay_202_0;
      shiftRegs_validIn_delay_204_0 <= shiftRegs_validIn_delay_203_0;
      shiftRegs_validIn_delay_205_0 <= shiftRegs_validIn_delay_204_0;
      shiftRegs_validIn_delay_206_0 <= shiftRegs_validIn_delay_205_0;
      shiftRegs_validIn_delay_207_0 <= shiftRegs_validIn_delay_206_0;
      shiftRegs_validIn_delay_208_0 <= shiftRegs_validIn_delay_207_0;
      shiftRegs_validIn_delay_209_0 <= shiftRegs_validIn_delay_208_0;
      shiftRegs_validIn_delay_210_0 <= shiftRegs_validIn_delay_209_0;
      shiftRegs_validIn_delay_211_0 <= shiftRegs_validIn_delay_210_0;
      shiftRegs_validIn_delay_212_0 <= shiftRegs_validIn_delay_211_0;
      shiftRegs_validIn_delay_213_0 <= shiftRegs_validIn_delay_212_0;
      shiftRegs_validIn_delay_214_0 <= shiftRegs_validIn_delay_213_0;
      shiftRegs_validIn_delay_215_0 <= shiftRegs_validIn_delay_214_0;
      shiftRegs_validIn_delay_216_0 <= shiftRegs_validIn_delay_215_0;
      shiftRegs_validIn_delay_217_0 <= shiftRegs_validIn_delay_216_0;
      shiftRegs_validIn_delay_218_0 <= shiftRegs_validIn_delay_217_0;
      shiftRegs_validIn_delay_219_0 <= shiftRegs_validIn_delay_218_0;
      shiftRegs_validIn_delay_220_0 <= shiftRegs_validIn_delay_219_0;
      shiftRegs_validIn_delay_221_0 <= shiftRegs_validIn_delay_220_0;
      shiftRegs_validIn_delay_222_0 <= shiftRegs_validIn_delay_221_0;
      shiftRegs_validIn_delay_223_0 <= shiftRegs_validIn_delay_222_0;
      shiftRegs_validIn_delay_224_0 <= shiftRegs_validIn_delay_223_0;
      shiftRegs_validIn_delay_225_0 <= shiftRegs_validIn_delay_224_0;
      shiftRegs_validIn_delay_226_0 <= shiftRegs_validIn_delay_225_0;
      shiftRegs_validIn_delay_227_0 <= shiftRegs_validIn_delay_226_0;
      shiftRegs_validIn_delay_228_0 <= shiftRegs_validIn_delay_227_0;
      shiftRegs_validIn_delay_229_0 <= shiftRegs_validIn_delay_228_0;
      shiftRegs_validIn_delay_230_0 <= shiftRegs_validIn_delay_229_0;
      shiftRegs_validIn_delay_231_0 <= shiftRegs_validIn_delay_230_0;
      shiftRegs_validIn_delay_232_0 <= shiftRegs_validIn_delay_231_0;
      shiftRegs_validIn_delay_233_0 <= shiftRegs_validIn_delay_232_0;
      shiftRegs_validIn_delay_234_0 <= shiftRegs_validIn_delay_233_0;
      shiftRegs_validIn_delay_235_0 <= shiftRegs_validIn_delay_234_0;
      shiftRegs_validIn_delay_236_0 <= shiftRegs_validIn_delay_235_0;
      shiftRegs_validIn_delay_237_0 <= shiftRegs_validIn_delay_236_0;
      shiftRegs_validIn_delay_238_0 <= shiftRegs_validIn_delay_237_0;
      shiftRegs_validIn_delay_239_0 <= shiftRegs_validIn_delay_238_0;
      shiftRegs_validIn_delay_240_0 <= shiftRegs_validIn_delay_239_0;
      shiftRegs_validIn_delay_241_0 <= shiftRegs_validIn_delay_240_0;
      shiftRegs_validIn_delay_242_0 <= shiftRegs_validIn_delay_241_0;
      shiftRegs_validIn_delay_243_0 <= shiftRegs_validIn_delay_242_0;
      shiftRegs_validIn_delay_244_0 <= shiftRegs_validIn_delay_243_0;
      shiftRegs_validIn_delay_245_0 <= shiftRegs_validIn_delay_244_0;
      shiftRegs_validIn_delay_246_0 <= shiftRegs_validIn_delay_245_0;
      shiftRegs_validIn_delay_247_0 <= shiftRegs_validIn_delay_246_0;
      shiftRegs_validIn_delay_248_0 <= shiftRegs_validIn_delay_247_0;
      shiftRegs_validIn_delay_249_0 <= shiftRegs_validIn_delay_248_0;
      shiftRegs_validIn_delay_250_0 <= shiftRegs_validIn_delay_249_0;
      shiftRegs_validIn_delay_251_0 <= shiftRegs_validIn_delay_250_0;
      shiftRegs_validIn_delay_252_0 <= shiftRegs_validIn_delay_251_0;
      shiftRegs_validIn_delay_253_0 <= shiftRegs_validIn_delay_252_0;
      shiftRegs_validIn_delay_254_0 <= shiftRegs_validIn_delay_253_0;
      shiftRegs_validOut_0 <= shiftRegs_validIn_delay_254_0;
      shiftRegs_validOut_delay_1_0 <= shiftRegs_validOut_0;
      shiftRegs_validOut_delay_2_0 <= shiftRegs_validOut_delay_1_0;
      shiftRegs_validOut_delay_3_0 <= shiftRegs_validOut_delay_2_0;
      shiftRegs_validOut_delay_4_0 <= shiftRegs_validOut_delay_3_0;
      shiftRegs_validOutFull_0 <= shiftRegs_validOut_delay_4_0;
      if(io_dataOut_ready) begin
        outputValid <= 1'b0;
      end
      flushing_flushCnt_value <= flushing_flushCnt_valueNext;
      flushing_flushCnt_willOverflowIfInc <= (flushing_flushCnt_valueNext == 17'h13fff);
      stage1_NCnt_value <= stage1_NCnt_valueNext;
      stage1_NCnt_willOverflowIfInc <= (stage1_NCnt_valueNext == 32'hffffffff);
      stage1_GCnt_value <= stage1_GCnt_valueNext;
      stage1_GCnt_willOverflowIfInc <= (stage1_GCnt_valueNext == 5'h13);
      stage1_emptyCnt_value <= stage1_emptyCnt_valueNext;
      stage1_emptyCnt_willOverflowIfInc <= (stage1_emptyCnt_valueNext == 9'h127);
      _zz_stage1_inputValid_0 <= (((((fsm_stateReg & fsm_enumDef_stage1) != 4'b0000) && (! stage1_waitReg)) && dataInBuffer_bufferOut_valid) && (_zz__zz_stage1_inputValid_0 != 13'h0));
      _zz_stage1_inputValid_0_1 <= _zz_stage1_inputValid_0;
      _zz_stage1_inputValid_0_2 <= _zz_stage1_inputValid_0_1;
      _zz_stage1_inputValid_0_3 <= _zz_stage1_inputValid_0_2;
      _zz_stage1_inputValid_0_4 <= _zz_stage1_inputValid_0_3;
      stage1_inputValid_0 <= _zz_stage1_inputValid_0_4;
      stage2_wCnt_value <= stage2_wCnt_valueNext;
      stage2_wCnt_willUnderflowIfDec <= (stage2_wCnt_valueNext == 12'h0);
      stage2_GCnt_value <= stage2_GCnt_valueNext;
      stage2_GCnt_willOverflowIfInc <= (stage2_GCnt_valueNext == 5'h13);
      stage2_calCnt_value <= stage2_calCnt_valueNext;
      stage2_calCnt_willUnderflowIfDec <= (stage2_calCnt_valueNext == 2'b00);
      stage2_waitCnt_value <= stage2_waitCnt_valueNext;
      stage2_waitCnt_willOverflowIfInc <= (stage2_waitCnt_valueNext == 9'h125);
      stage3_GCnt_value <= stage3_GCnt_valueNext;
      stage3_GCnt_willUnderflowIfDec <= (stage3_GCnt_valueNext == 5'h01);
      stage3_doubleCnt_value <= stage3_doubleCnt_valueNext;
      stage3_doubleCnt_willOverflowIfInc <= (stage3_doubleCnt_valueNext == 4'b1100);
      stage3_doubleWaitCnt_value <= stage3_doubleWaitCnt_valueNext;
      stage3_doubleWaitCnt_willOverflowIfInc <= (stage3_doubleWaitCnt_valueNext == 9'h127);
      stage3_addWaitCnt_value <= stage3_addWaitCnt_valueNext;
      stage3_addWaitCnt_willOverflowIfInc <= (stage3_addWaitCnt_valueNext == 9'h127);
      fsm_stateReg <= fsm_stateNext;
      (* parallel_case *)
      case(1) // synthesis parallel_case
        (((fsm_stateReg) & fsm_enumDef_stage1) == fsm_enumDef_stage1) : begin
          if(when_Pippenger_l153) begin
            if(dataInBuffer_bufferOut_valid) begin
              if(stage1_GCnt_willOverflowIfInc) begin
                if(dataInBuffer_bufferOut_payload_last) begin
                  stage1_waitReg <= 1'b1;
                end
              end
              stage1_needAdd1_0 <= (|stage1_inputBarrelID_0[13 : 12]);
            end
          end else begin
            if(!when_Pippenger_l168) begin
              if(stage1_emptyCnt_willOverflowIfInc) begin
                stage1_waitReg <= 1'b0;
              end
            end
          end
        end
        (((fsm_stateReg) & fsm_enumDef_stage2) == fsm_enumDef_stage2) : begin
          if(when_Pippenger_l207) begin
            if(stage2_calCnt_willUnderflowIfDec) begin
              if(stage2_GCnt_willOverflowIfInc) begin
                stage2_waitReg <= 1'b1;
              end
            end
          end else begin
            if(stage2_waitCnt_willOverflowIfInc) begin
              stage2_waitReg <= 1'b0;
            end
          end
        end
        (((fsm_stateReg) & fsm_enumDef_stage3) == fsm_enumDef_stage3) : begin
          if(when_Pippenger_l249) begin
            if(stage3_doubleWaitCnt_willOverflowIfInc) begin
              if(stage3_doubleCnt_willOverflowIfInc) begin
                stage3_addReg <= 1'b1;
              end
            end
          end else begin
            if(stage3_addWaitCnt_willOverflowIfInc) begin
              stage3_addReg <= 1'b0;
              if(stage3_GCnt_willUnderflowIfDec) begin
                outputValid <= 1'b1;
              end
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if(io_dataIn_ready) begin
      dataInBuffer_dataReg_last <= io_dataIn_payload_last;
      dataInBuffer_dataReg_fragment_P_X <= io_dataIn_payload_fragment_P_X;
      dataInBuffer_dataReg_fragment_P_Y <= io_dataIn_payload_fragment_P_Y;
      dataInBuffer_dataReg_fragment_P_Z <= io_dataIn_payload_fragment_P_Z;
      dataInBuffer_dataReg_fragment_P_T <= io_dataIn_payload_fragment_P_T;
      dataInBuffer_dataReg_fragment_K <= io_dataIn_payload_fragment_K;
    end else begin
      if(dataInBuffer_shift) begin
        dataInBuffer_dataReg_fragment_K <= {13'd0, _zz_dataInBuffer_dataReg_fragment_K};
      end
    end
    shiftRegs_addressIn_delay_1_0 <= shiftRegs_addressIn_0;
    shiftRegs_addressIn_delay_2_0 <= shiftRegs_addressIn_delay_1_0;
    shiftRegs_addressIn_delay_3_0 <= shiftRegs_addressIn_delay_2_0;
    shiftRegs_addressIn_delay_4_0 <= shiftRegs_addressIn_delay_3_0;
    shiftRegs_addressIn_delay_5_0 <= shiftRegs_addressIn_delay_4_0;
    shiftRegs_addressIn_delay_6_0 <= shiftRegs_addressIn_delay_5_0;
    shiftRegs_addressIn_delay_7_0 <= shiftRegs_addressIn_delay_6_0;
    shiftRegs_addressIn_delay_8_0 <= shiftRegs_addressIn_delay_7_0;
    shiftRegs_addressIn_delay_9_0 <= shiftRegs_addressIn_delay_8_0;
    shiftRegs_addressIn_delay_10_0 <= shiftRegs_addressIn_delay_9_0;
    shiftRegs_addressIn_delay_11_0 <= shiftRegs_addressIn_delay_10_0;
    shiftRegs_addressIn_delay_12_0 <= shiftRegs_addressIn_delay_11_0;
    shiftRegs_addressIn_delay_13_0 <= shiftRegs_addressIn_delay_12_0;
    shiftRegs_addressIn_delay_14_0 <= shiftRegs_addressIn_delay_13_0;
    shiftRegs_addressIn_delay_15_0 <= shiftRegs_addressIn_delay_14_0;
    shiftRegs_addressIn_delay_16_0 <= shiftRegs_addressIn_delay_15_0;
    shiftRegs_addressIn_delay_17_0 <= shiftRegs_addressIn_delay_16_0;
    shiftRegs_addressIn_delay_18_0 <= shiftRegs_addressIn_delay_17_0;
    shiftRegs_addressIn_delay_19_0 <= shiftRegs_addressIn_delay_18_0;
    shiftRegs_addressIn_delay_20_0 <= shiftRegs_addressIn_delay_19_0;
    shiftRegs_addressIn_delay_21_0 <= shiftRegs_addressIn_delay_20_0;
    shiftRegs_addressIn_delay_22_0 <= shiftRegs_addressIn_delay_21_0;
    shiftRegs_addressIn_delay_23_0 <= shiftRegs_addressIn_delay_22_0;
    shiftRegs_addressIn_delay_24_0 <= shiftRegs_addressIn_delay_23_0;
    shiftRegs_addressIn_delay_25_0 <= shiftRegs_addressIn_delay_24_0;
    shiftRegs_addressIn_delay_26_0 <= shiftRegs_addressIn_delay_25_0;
    shiftRegs_addressIn_delay_27_0 <= shiftRegs_addressIn_delay_26_0;
    shiftRegs_addressIn_delay_28_0 <= shiftRegs_addressIn_delay_27_0;
    shiftRegs_addressIn_delay_29_0 <= shiftRegs_addressIn_delay_28_0;
    shiftRegs_addressIn_delay_30_0 <= shiftRegs_addressIn_delay_29_0;
    shiftRegs_addressIn_delay_31_0 <= shiftRegs_addressIn_delay_30_0;
    shiftRegs_addressIn_delay_32_0 <= shiftRegs_addressIn_delay_31_0;
    shiftRegs_addressIn_delay_33_0 <= shiftRegs_addressIn_delay_32_0;
    shiftRegs_addressIn_delay_34_0 <= shiftRegs_addressIn_delay_33_0;
    shiftRegs_addressIn_delay_35_0 <= shiftRegs_addressIn_delay_34_0;
    shiftRegs_addressIn_delay_36_0 <= shiftRegs_addressIn_delay_35_0;
    shiftRegs_addressIn_delay_37_0 <= shiftRegs_addressIn_delay_36_0;
    shiftRegs_addressIn_delay_38_0 <= shiftRegs_addressIn_delay_37_0;
    shiftRegs_addressIn_delay_39_0 <= shiftRegs_addressIn_delay_38_0;
    shiftRegs_addressIn_delay_40_0 <= shiftRegs_addressIn_delay_39_0;
    shiftRegs_addressIn_delay_41_0 <= shiftRegs_addressIn_delay_40_0;
    shiftRegs_addressIn_delay_42_0 <= shiftRegs_addressIn_delay_41_0;
    shiftRegs_addressIn_delay_43_0 <= shiftRegs_addressIn_delay_42_0;
    shiftRegs_addressIn_delay_44_0 <= shiftRegs_addressIn_delay_43_0;
    shiftRegs_addressIn_delay_45_0 <= shiftRegs_addressIn_delay_44_0;
    shiftRegs_addressIn_delay_46_0 <= shiftRegs_addressIn_delay_45_0;
    shiftRegs_addressIn_delay_47_0 <= shiftRegs_addressIn_delay_46_0;
    shiftRegs_addressIn_delay_48_0 <= shiftRegs_addressIn_delay_47_0;
    shiftRegs_addressIn_delay_49_0 <= shiftRegs_addressIn_delay_48_0;
    shiftRegs_addressIn_delay_50_0 <= shiftRegs_addressIn_delay_49_0;
    shiftRegs_addressIn_delay_51_0 <= shiftRegs_addressIn_delay_50_0;
    shiftRegs_addressIn_delay_52_0 <= shiftRegs_addressIn_delay_51_0;
    shiftRegs_addressIn_delay_53_0 <= shiftRegs_addressIn_delay_52_0;
    shiftRegs_addressIn_delay_54_0 <= shiftRegs_addressIn_delay_53_0;
    shiftRegs_addressIn_delay_55_0 <= shiftRegs_addressIn_delay_54_0;
    shiftRegs_addressIn_delay_56_0 <= shiftRegs_addressIn_delay_55_0;
    shiftRegs_addressIn_delay_57_0 <= shiftRegs_addressIn_delay_56_0;
    shiftRegs_addressIn_delay_58_0 <= shiftRegs_addressIn_delay_57_0;
    shiftRegs_addressIn_delay_59_0 <= shiftRegs_addressIn_delay_58_0;
    shiftRegs_addressIn_delay_60_0 <= shiftRegs_addressIn_delay_59_0;
    shiftRegs_addressIn_delay_61_0 <= shiftRegs_addressIn_delay_60_0;
    shiftRegs_addressIn_delay_62_0 <= shiftRegs_addressIn_delay_61_0;
    shiftRegs_addressIn_delay_63_0 <= shiftRegs_addressIn_delay_62_0;
    shiftRegs_addressIn_delay_64_0 <= shiftRegs_addressIn_delay_63_0;
    shiftRegs_addressIn_delay_65_0 <= shiftRegs_addressIn_delay_64_0;
    shiftRegs_addressIn_delay_66_0 <= shiftRegs_addressIn_delay_65_0;
    shiftRegs_addressIn_delay_67_0 <= shiftRegs_addressIn_delay_66_0;
    shiftRegs_addressIn_delay_68_0 <= shiftRegs_addressIn_delay_67_0;
    shiftRegs_addressIn_delay_69_0 <= shiftRegs_addressIn_delay_68_0;
    shiftRegs_addressIn_delay_70_0 <= shiftRegs_addressIn_delay_69_0;
    shiftRegs_addressIn_delay_71_0 <= shiftRegs_addressIn_delay_70_0;
    shiftRegs_addressIn_delay_72_0 <= shiftRegs_addressIn_delay_71_0;
    shiftRegs_addressIn_delay_73_0 <= shiftRegs_addressIn_delay_72_0;
    shiftRegs_addressIn_delay_74_0 <= shiftRegs_addressIn_delay_73_0;
    shiftRegs_addressIn_delay_75_0 <= shiftRegs_addressIn_delay_74_0;
    shiftRegs_addressIn_delay_76_0 <= shiftRegs_addressIn_delay_75_0;
    shiftRegs_addressIn_delay_77_0 <= shiftRegs_addressIn_delay_76_0;
    shiftRegs_addressIn_delay_78_0 <= shiftRegs_addressIn_delay_77_0;
    shiftRegs_addressIn_delay_79_0 <= shiftRegs_addressIn_delay_78_0;
    shiftRegs_addressIn_delay_80_0 <= shiftRegs_addressIn_delay_79_0;
    shiftRegs_addressIn_delay_81_0 <= shiftRegs_addressIn_delay_80_0;
    shiftRegs_addressIn_delay_82_0 <= shiftRegs_addressIn_delay_81_0;
    shiftRegs_addressIn_delay_83_0 <= shiftRegs_addressIn_delay_82_0;
    shiftRegs_addressIn_delay_84_0 <= shiftRegs_addressIn_delay_83_0;
    shiftRegs_addressIn_delay_85_0 <= shiftRegs_addressIn_delay_84_0;
    shiftRegs_addressIn_delay_86_0 <= shiftRegs_addressIn_delay_85_0;
    shiftRegs_addressIn_delay_87_0 <= shiftRegs_addressIn_delay_86_0;
    shiftRegs_addressIn_delay_88_0 <= shiftRegs_addressIn_delay_87_0;
    shiftRegs_addressIn_delay_89_0 <= shiftRegs_addressIn_delay_88_0;
    shiftRegs_addressIn_delay_90_0 <= shiftRegs_addressIn_delay_89_0;
    shiftRegs_addressIn_delay_91_0 <= shiftRegs_addressIn_delay_90_0;
    shiftRegs_addressIn_delay_92_0 <= shiftRegs_addressIn_delay_91_0;
    shiftRegs_addressIn_delay_93_0 <= shiftRegs_addressIn_delay_92_0;
    shiftRegs_addressIn_delay_94_0 <= shiftRegs_addressIn_delay_93_0;
    shiftRegs_addressIn_delay_95_0 <= shiftRegs_addressIn_delay_94_0;
    shiftRegs_addressIn_delay_96_0 <= shiftRegs_addressIn_delay_95_0;
    shiftRegs_addressIn_delay_97_0 <= shiftRegs_addressIn_delay_96_0;
    shiftRegs_addressIn_delay_98_0 <= shiftRegs_addressIn_delay_97_0;
    shiftRegs_addressIn_delay_99_0 <= shiftRegs_addressIn_delay_98_0;
    shiftRegs_addressIn_delay_100_0 <= shiftRegs_addressIn_delay_99_0;
    shiftRegs_addressIn_delay_101_0 <= shiftRegs_addressIn_delay_100_0;
    shiftRegs_addressIn_delay_102_0 <= shiftRegs_addressIn_delay_101_0;
    shiftRegs_addressIn_delay_103_0 <= shiftRegs_addressIn_delay_102_0;
    shiftRegs_addressIn_delay_104_0 <= shiftRegs_addressIn_delay_103_0;
    shiftRegs_addressIn_delay_105_0 <= shiftRegs_addressIn_delay_104_0;
    shiftRegs_addressIn_delay_106_0 <= shiftRegs_addressIn_delay_105_0;
    shiftRegs_addressIn_delay_107_0 <= shiftRegs_addressIn_delay_106_0;
    shiftRegs_addressIn_delay_108_0 <= shiftRegs_addressIn_delay_107_0;
    shiftRegs_addressIn_delay_109_0 <= shiftRegs_addressIn_delay_108_0;
    shiftRegs_addressIn_delay_110_0 <= shiftRegs_addressIn_delay_109_0;
    shiftRegs_addressIn_delay_111_0 <= shiftRegs_addressIn_delay_110_0;
    shiftRegs_addressIn_delay_112_0 <= shiftRegs_addressIn_delay_111_0;
    shiftRegs_addressIn_delay_113_0 <= shiftRegs_addressIn_delay_112_0;
    shiftRegs_addressIn_delay_114_0 <= shiftRegs_addressIn_delay_113_0;
    shiftRegs_addressIn_delay_115_0 <= shiftRegs_addressIn_delay_114_0;
    shiftRegs_addressIn_delay_116_0 <= shiftRegs_addressIn_delay_115_0;
    shiftRegs_addressIn_delay_117_0 <= shiftRegs_addressIn_delay_116_0;
    shiftRegs_addressIn_delay_118_0 <= shiftRegs_addressIn_delay_117_0;
    shiftRegs_addressIn_delay_119_0 <= shiftRegs_addressIn_delay_118_0;
    shiftRegs_addressIn_delay_120_0 <= shiftRegs_addressIn_delay_119_0;
    shiftRegs_addressIn_delay_121_0 <= shiftRegs_addressIn_delay_120_0;
    shiftRegs_addressIn_delay_122_0 <= shiftRegs_addressIn_delay_121_0;
    shiftRegs_addressIn_delay_123_0 <= shiftRegs_addressIn_delay_122_0;
    shiftRegs_addressIn_delay_124_0 <= shiftRegs_addressIn_delay_123_0;
    shiftRegs_addressIn_delay_125_0 <= shiftRegs_addressIn_delay_124_0;
    shiftRegs_addressIn_delay_126_0 <= shiftRegs_addressIn_delay_125_0;
    shiftRegs_addressIn_delay_127_0 <= shiftRegs_addressIn_delay_126_0;
    shiftRegs_addressIn_delay_128_0 <= shiftRegs_addressIn_delay_127_0;
    shiftRegs_addressIn_delay_129_0 <= shiftRegs_addressIn_delay_128_0;
    shiftRegs_addressIn_delay_130_0 <= shiftRegs_addressIn_delay_129_0;
    shiftRegs_addressIn_delay_131_0 <= shiftRegs_addressIn_delay_130_0;
    shiftRegs_addressIn_delay_132_0 <= shiftRegs_addressIn_delay_131_0;
    shiftRegs_addressIn_delay_133_0 <= shiftRegs_addressIn_delay_132_0;
    shiftRegs_addressIn_delay_134_0 <= shiftRegs_addressIn_delay_133_0;
    shiftRegs_addressIn_delay_135_0 <= shiftRegs_addressIn_delay_134_0;
    shiftRegs_addressIn_delay_136_0 <= shiftRegs_addressIn_delay_135_0;
    shiftRegs_addressIn_delay_137_0 <= shiftRegs_addressIn_delay_136_0;
    shiftRegs_addressIn_delay_138_0 <= shiftRegs_addressIn_delay_137_0;
    shiftRegs_addressIn_delay_139_0 <= shiftRegs_addressIn_delay_138_0;
    shiftRegs_addressIn_delay_140_0 <= shiftRegs_addressIn_delay_139_0;
    shiftRegs_addressIn_delay_141_0 <= shiftRegs_addressIn_delay_140_0;
    shiftRegs_addressIn_delay_142_0 <= shiftRegs_addressIn_delay_141_0;
    shiftRegs_addressIn_delay_143_0 <= shiftRegs_addressIn_delay_142_0;
    shiftRegs_addressIn_delay_144_0 <= shiftRegs_addressIn_delay_143_0;
    shiftRegs_addressIn_delay_145_0 <= shiftRegs_addressIn_delay_144_0;
    shiftRegs_addressIn_delay_146_0 <= shiftRegs_addressIn_delay_145_0;
    shiftRegs_addressIn_delay_147_0 <= shiftRegs_addressIn_delay_146_0;
    shiftRegs_addressIn_delay_148_0 <= shiftRegs_addressIn_delay_147_0;
    shiftRegs_addressIn_delay_149_0 <= shiftRegs_addressIn_delay_148_0;
    shiftRegs_addressIn_delay_150_0 <= shiftRegs_addressIn_delay_149_0;
    shiftRegs_addressIn_delay_151_0 <= shiftRegs_addressIn_delay_150_0;
    shiftRegs_addressIn_delay_152_0 <= shiftRegs_addressIn_delay_151_0;
    shiftRegs_addressIn_delay_153_0 <= shiftRegs_addressIn_delay_152_0;
    shiftRegs_addressIn_delay_154_0 <= shiftRegs_addressIn_delay_153_0;
    shiftRegs_addressIn_delay_155_0 <= shiftRegs_addressIn_delay_154_0;
    shiftRegs_addressIn_delay_156_0 <= shiftRegs_addressIn_delay_155_0;
    shiftRegs_addressIn_delay_157_0 <= shiftRegs_addressIn_delay_156_0;
    shiftRegs_addressIn_delay_158_0 <= shiftRegs_addressIn_delay_157_0;
    shiftRegs_addressIn_delay_159_0 <= shiftRegs_addressIn_delay_158_0;
    shiftRegs_addressIn_delay_160_0 <= shiftRegs_addressIn_delay_159_0;
    shiftRegs_addressIn_delay_161_0 <= shiftRegs_addressIn_delay_160_0;
    shiftRegs_addressIn_delay_162_0 <= shiftRegs_addressIn_delay_161_0;
    shiftRegs_addressIn_delay_163_0 <= shiftRegs_addressIn_delay_162_0;
    shiftRegs_addressIn_delay_164_0 <= shiftRegs_addressIn_delay_163_0;
    shiftRegs_addressIn_delay_165_0 <= shiftRegs_addressIn_delay_164_0;
    shiftRegs_addressIn_delay_166_0 <= shiftRegs_addressIn_delay_165_0;
    shiftRegs_addressIn_delay_167_0 <= shiftRegs_addressIn_delay_166_0;
    shiftRegs_addressIn_delay_168_0 <= shiftRegs_addressIn_delay_167_0;
    shiftRegs_addressIn_delay_169_0 <= shiftRegs_addressIn_delay_168_0;
    shiftRegs_addressIn_delay_170_0 <= shiftRegs_addressIn_delay_169_0;
    shiftRegs_addressIn_delay_171_0 <= shiftRegs_addressIn_delay_170_0;
    shiftRegs_addressIn_delay_172_0 <= shiftRegs_addressIn_delay_171_0;
    shiftRegs_addressIn_delay_173_0 <= shiftRegs_addressIn_delay_172_0;
    shiftRegs_addressIn_delay_174_0 <= shiftRegs_addressIn_delay_173_0;
    shiftRegs_addressIn_delay_175_0 <= shiftRegs_addressIn_delay_174_0;
    shiftRegs_addressIn_delay_176_0 <= shiftRegs_addressIn_delay_175_0;
    shiftRegs_addressIn_delay_177_0 <= shiftRegs_addressIn_delay_176_0;
    shiftRegs_addressIn_delay_178_0 <= shiftRegs_addressIn_delay_177_0;
    shiftRegs_addressIn_delay_179_0 <= shiftRegs_addressIn_delay_178_0;
    shiftRegs_addressIn_delay_180_0 <= shiftRegs_addressIn_delay_179_0;
    shiftRegs_addressIn_delay_181_0 <= shiftRegs_addressIn_delay_180_0;
    shiftRegs_addressIn_delay_182_0 <= shiftRegs_addressIn_delay_181_0;
    shiftRegs_addressIn_delay_183_0 <= shiftRegs_addressIn_delay_182_0;
    shiftRegs_addressIn_delay_184_0 <= shiftRegs_addressIn_delay_183_0;
    shiftRegs_addressIn_delay_185_0 <= shiftRegs_addressIn_delay_184_0;
    shiftRegs_addressIn_delay_186_0 <= shiftRegs_addressIn_delay_185_0;
    shiftRegs_addressIn_delay_187_0 <= shiftRegs_addressIn_delay_186_0;
    shiftRegs_addressIn_delay_188_0 <= shiftRegs_addressIn_delay_187_0;
    shiftRegs_addressIn_delay_189_0 <= shiftRegs_addressIn_delay_188_0;
    shiftRegs_addressIn_delay_190_0 <= shiftRegs_addressIn_delay_189_0;
    shiftRegs_addressIn_delay_191_0 <= shiftRegs_addressIn_delay_190_0;
    shiftRegs_addressIn_delay_192_0 <= shiftRegs_addressIn_delay_191_0;
    shiftRegs_addressIn_delay_193_0 <= shiftRegs_addressIn_delay_192_0;
    shiftRegs_addressIn_delay_194_0 <= shiftRegs_addressIn_delay_193_0;
    shiftRegs_addressIn_delay_195_0 <= shiftRegs_addressIn_delay_194_0;
    shiftRegs_addressIn_delay_196_0 <= shiftRegs_addressIn_delay_195_0;
    shiftRegs_addressIn_delay_197_0 <= shiftRegs_addressIn_delay_196_0;
    shiftRegs_addressIn_delay_198_0 <= shiftRegs_addressIn_delay_197_0;
    shiftRegs_addressIn_delay_199_0 <= shiftRegs_addressIn_delay_198_0;
    shiftRegs_addressIn_delay_200_0 <= shiftRegs_addressIn_delay_199_0;
    shiftRegs_addressIn_delay_201_0 <= shiftRegs_addressIn_delay_200_0;
    shiftRegs_addressIn_delay_202_0 <= shiftRegs_addressIn_delay_201_0;
    shiftRegs_addressIn_delay_203_0 <= shiftRegs_addressIn_delay_202_0;
    shiftRegs_addressIn_delay_204_0 <= shiftRegs_addressIn_delay_203_0;
    shiftRegs_addressIn_delay_205_0 <= shiftRegs_addressIn_delay_204_0;
    shiftRegs_addressIn_delay_206_0 <= shiftRegs_addressIn_delay_205_0;
    shiftRegs_addressIn_delay_207_0 <= shiftRegs_addressIn_delay_206_0;
    shiftRegs_addressIn_delay_208_0 <= shiftRegs_addressIn_delay_207_0;
    shiftRegs_addressIn_delay_209_0 <= shiftRegs_addressIn_delay_208_0;
    shiftRegs_addressIn_delay_210_0 <= shiftRegs_addressIn_delay_209_0;
    shiftRegs_addressIn_delay_211_0 <= shiftRegs_addressIn_delay_210_0;
    shiftRegs_addressIn_delay_212_0 <= shiftRegs_addressIn_delay_211_0;
    shiftRegs_addressIn_delay_213_0 <= shiftRegs_addressIn_delay_212_0;
    shiftRegs_addressIn_delay_214_0 <= shiftRegs_addressIn_delay_213_0;
    shiftRegs_addressIn_delay_215_0 <= shiftRegs_addressIn_delay_214_0;
    shiftRegs_addressIn_delay_216_0 <= shiftRegs_addressIn_delay_215_0;
    shiftRegs_addressIn_delay_217_0 <= shiftRegs_addressIn_delay_216_0;
    shiftRegs_addressIn_delay_218_0 <= shiftRegs_addressIn_delay_217_0;
    shiftRegs_addressIn_delay_219_0 <= shiftRegs_addressIn_delay_218_0;
    shiftRegs_addressIn_delay_220_0 <= shiftRegs_addressIn_delay_219_0;
    shiftRegs_addressIn_delay_221_0 <= shiftRegs_addressIn_delay_220_0;
    shiftRegs_addressIn_delay_222_0 <= shiftRegs_addressIn_delay_221_0;
    shiftRegs_addressIn_delay_223_0 <= shiftRegs_addressIn_delay_222_0;
    shiftRegs_addressIn_delay_224_0 <= shiftRegs_addressIn_delay_223_0;
    shiftRegs_addressIn_delay_225_0 <= shiftRegs_addressIn_delay_224_0;
    shiftRegs_addressIn_delay_226_0 <= shiftRegs_addressIn_delay_225_0;
    shiftRegs_addressIn_delay_227_0 <= shiftRegs_addressIn_delay_226_0;
    shiftRegs_addressIn_delay_228_0 <= shiftRegs_addressIn_delay_227_0;
    shiftRegs_addressIn_delay_229_0 <= shiftRegs_addressIn_delay_228_0;
    shiftRegs_addressIn_delay_230_0 <= shiftRegs_addressIn_delay_229_0;
    shiftRegs_addressIn_delay_231_0 <= shiftRegs_addressIn_delay_230_0;
    shiftRegs_addressIn_delay_232_0 <= shiftRegs_addressIn_delay_231_0;
    shiftRegs_addressIn_delay_233_0 <= shiftRegs_addressIn_delay_232_0;
    shiftRegs_addressIn_delay_234_0 <= shiftRegs_addressIn_delay_233_0;
    shiftRegs_addressIn_delay_235_0 <= shiftRegs_addressIn_delay_234_0;
    shiftRegs_addressIn_delay_236_0 <= shiftRegs_addressIn_delay_235_0;
    shiftRegs_addressIn_delay_237_0 <= shiftRegs_addressIn_delay_236_0;
    shiftRegs_addressIn_delay_238_0 <= shiftRegs_addressIn_delay_237_0;
    shiftRegs_addressIn_delay_239_0 <= shiftRegs_addressIn_delay_238_0;
    shiftRegs_addressIn_delay_240_0 <= shiftRegs_addressIn_delay_239_0;
    shiftRegs_addressIn_delay_241_0 <= shiftRegs_addressIn_delay_240_0;
    shiftRegs_addressIn_delay_242_0 <= shiftRegs_addressIn_delay_241_0;
    shiftRegs_addressIn_delay_243_0 <= shiftRegs_addressIn_delay_242_0;
    shiftRegs_addressIn_delay_244_0 <= shiftRegs_addressIn_delay_243_0;
    shiftRegs_addressIn_delay_245_0 <= shiftRegs_addressIn_delay_244_0;
    shiftRegs_addressIn_delay_246_0 <= shiftRegs_addressIn_delay_245_0;
    shiftRegs_addressIn_delay_247_0 <= shiftRegs_addressIn_delay_246_0;
    shiftRegs_addressIn_delay_248_0 <= shiftRegs_addressIn_delay_247_0;
    shiftRegs_addressIn_delay_249_0 <= shiftRegs_addressIn_delay_248_0;
    shiftRegs_addressIn_delay_250_0 <= shiftRegs_addressIn_delay_249_0;
    shiftRegs_addressIn_delay_251_0 <= shiftRegs_addressIn_delay_250_0;
    shiftRegs_addressIn_delay_252_0 <= shiftRegs_addressIn_delay_251_0;
    shiftRegs_addressIn_delay_253_0 <= shiftRegs_addressIn_delay_252_0;
    shiftRegs_addressIn_delay_254_0 <= shiftRegs_addressIn_delay_253_0;
    shiftRegs_addressOut_0 <= shiftRegs_addressIn_delay_254_0;
    shiftRegs_addressOut_delay_1_0 <= shiftRegs_addressOut_0;
    shiftRegs_addressOut_delay_2_0 <= shiftRegs_addressOut_delay_1_0;
    shiftRegs_addressOut_delay_3_0 <= shiftRegs_addressOut_delay_2_0;
    shiftRegs_addressOut_delay_4_0 <= shiftRegs_addressOut_delay_3_0;
    shiftRegs_addressOutFull_0 <= shiftRegs_addressOut_delay_4_0;
    pAddPort_0_s_regNext_X <= pAddPort_0_s_X;
    pAddPort_0_s_regNext_Y <= pAddPort_0_s_Y;
    pAddPort_0_s_regNext_Z <= pAddPort_0_s_Z;
    pAddPort_0_s_regNext_T <= pAddPort_0_s_T;
    _zz_stage1_inputAddress_0 <= {stage1_GCnt_value,stage1_inputBarrelIDAbs_0};
    _zz_stage1_inputAddress_0_1 <= _zz_stage1_inputAddress_0;
    _zz_stage1_inputAddress_0_2 <= _zz_stage1_inputAddress_0_1;
    _zz_stage1_inputAddress_0_3 <= _zz_stage1_inputAddress_0_2;
    _zz_stage1_inputAddress_0_4 <= _zz_stage1_inputAddress_0_3;
    stage1_inputAddress_0 <= _zz_stage1_inputAddress_0_4;
    _zz_stage1_inputData_0_X <= stage1_inputBarrelID_0[12];
    _zz_stage1_inputData_0_X_1 <= _zz_stage1_inputData_0_X;
    _zz_stage1_inputData_0_X_2 <= _zz_stage1_inputData_0_X_1;
    _zz_stage1_inputData_0_X_3 <= _zz_stage1_inputData_0_X_2;
    _zz_stage1_inputData_0_X_4 <= _zz_stage1_inputData_0_X_3;
    _zz_stage1_inputData_0_X_5 <= _zz_stage1_inputData_0_X_4;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_X <= dataInBuffer_bufferOut_payload_fragment_P_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y <= dataInBuffer_bufferOut_payload_fragment_P_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z <= dataInBuffer_bufferOut_payload_fragment_P_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_1_T <= dataInBuffer_bufferOut_payload_fragment_P_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_2_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_1_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_3_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_2_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_4_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_3_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_5_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_4_T;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_X <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_X;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_Y <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_Y;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_Z <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_Z;
    dataInBuffer_bufferOut_payload_fragment_P_delay_6_T <= dataInBuffer_bufferOut_payload_fragment_P_delay_5_T;
  end

  always @(posedge clk) begin
    stage1_inputValid_0_delay_1 <= stage1_inputValid_0;
    stage1_inputValid_0_delay_2 <= stage1_inputValid_0_delay_1;
    stage1_inputValid_0_delay_3 <= stage1_inputValid_0_delay_2;
    stage1_inputValid_0_delay_4 <= stage1_inputValid_0_delay_3;
    stage1_inputValid_0_delay_5 <= stage1_inputValid_0_delay_4;
    stage1_inputAddress_0_delay_1 <= stage1_inputAddress_0;
    stage1_inputAddress_0_delay_2 <= stage1_inputAddress_0_delay_1;
    stage1_inputAddress_0_delay_3 <= stage1_inputAddress_0_delay_2;
    stage1_inputAddress_0_delay_4 <= stage1_inputAddress_0_delay_3;
    stage1_inputAddress_0_delay_5 <= stage1_inputAddress_0_delay_4;
    stage1_inputData_0_delay_1_X <= stage1_inputData_0_X;
    stage1_inputData_0_delay_1_Y <= stage1_inputData_0_Y;
    stage1_inputData_0_delay_1_Z <= stage1_inputData_0_Z;
    stage1_inputData_0_delay_1_T <= stage1_inputData_0_T;
    stage1_inputData_0_delay_2_X <= stage1_inputData_0_delay_1_X;
    stage1_inputData_0_delay_2_Y <= stage1_inputData_0_delay_1_Y;
    stage1_inputData_0_delay_2_Z <= stage1_inputData_0_delay_1_Z;
    stage1_inputData_0_delay_2_T <= stage1_inputData_0_delay_1_T;
    stage1_inputData_0_delay_3_X <= stage1_inputData_0_delay_2_X;
    stage1_inputData_0_delay_3_Y <= stage1_inputData_0_delay_2_Y;
    stage1_inputData_0_delay_3_Z <= stage1_inputData_0_delay_2_Z;
    stage1_inputData_0_delay_3_T <= stage1_inputData_0_delay_2_T;
    stage1_inputData_0_delay_4_X <= stage1_inputData_0_delay_3_X;
    stage1_inputData_0_delay_4_Y <= stage1_inputData_0_delay_3_Y;
    stage1_inputData_0_delay_4_Z <= stage1_inputData_0_delay_3_Z;
    stage1_inputData_0_delay_4_T <= stage1_inputData_0_delay_3_T;
    stage1_inputData_0_delay_5_X <= stage1_inputData_0_delay_4_X;
    stage1_inputData_0_delay_5_Y <= stage1_inputData_0_delay_4_Y;
    stage1_inputData_0_delay_5_Z <= stage1_inputData_0_delay_4_Z;
    stage1_inputData_0_delay_5_T <= stage1_inputData_0_delay_4_T;
    _zz_io_dataIn_0_valid <= (stage1_inputValid_0 && (stage1_inputAddress_0 == shiftRegs_addressOut_0));
    _zz_io_dataIn_0_valid_1 <= _zz_io_dataIn_0_valid;
    _zz_io_dataIn_0_valid_2 <= _zz_io_dataIn_0_valid_1;
    _zz_io_dataIn_0_valid_3 <= _zz_io_dataIn_0_valid_2;
    _zz_io_dataIn_0_valid_4 <= _zz_io_dataIn_0_valid_3;
    _zz_io_dataIn_0_payload_a_X <= (stage1_inputValid_0 && (stage1_inputAddress_0 == shiftRegs_addressOut_0));
    _zz_io_dataIn_0_payload_a_X_1 <= _zz_io_dataIn_0_payload_a_X;
    _zz_io_dataIn_0_payload_a_X_2 <= _zz_io_dataIn_0_payload_a_X_1;
    _zz_io_dataIn_0_payload_a_X_3 <= _zz_io_dataIn_0_payload_a_X_2;
    _zz_io_dataIn_0_payload_a_X_4 <= _zz_io_dataIn_0_payload_a_X_3;
    _zz_io_dataIn_0_payload_a_X_5 <= _zz_io_dataIn_0_payload_a_X_4;
    _zz_io_dataIn_0_payload_a_X_6 <= _zz_io_dataIn_0_payload_a_X_5;
    _zz_io_dataIn_0_payload_a_X_7 <= _zz_io_dataIn_0_payload_a_X_6;
    _zz_io_dataIn_0_payload_a_X_8 <= _zz_io_dataIn_0_payload_a_X_7;
    _zz_io_dataIn_0_payload_a_X_9 <= _zz_io_dataIn_0_payload_a_X_8;
    _zz_io_dataIn_0_payload_a_X_10 <= _zz_io_dataIn_0_payload_a_X_9;
    _zz_io_dataIn_0_payload_a_X_11 <= _zz_io_dataIn_0_payload_a_X_10;
    _zz_io_dataIn_0_payload_a_X_12 <= _zz_io_dataIn_0_payload_a_X_11;
    _zz_io_dataIn_0_payload_a_X_13 <= _zz_io_dataIn_0_payload_a_X_12;
    _zz_io_dataIn_0_payload_a_X_14 <= _zz_io_dataIn_0_payload_a_X_13;
    _zz_io_dataIn_0_payload_a_X_15 <= _zz_io_dataIn_0_payload_a_X_14;
    _zz_io_dataIn_0_payload_a_X_16 <= _zz_io_dataIn_0_payload_a_X_15;
    _zz_io_dataIn_0_payload_a_X_17 <= _zz_io_dataIn_0_payload_a_X_16;
    _zz_io_dataIn_0_payload_a_X_18 <= _zz_io_dataIn_0_payload_a_X_17;
    _zz_io_dataIn_0_payload_a_X_19 <= _zz_io_dataIn_0_payload_a_X_18;
    _zz_io_dataIn_0_payload_a_X_20 <= _zz_io_dataIn_0_payload_a_X_19;
    _zz_io_dataIn_0_payload_a_X_21 <= _zz_io_dataIn_0_payload_a_X_20;
    _zz_io_dataIn_0_payload_a_X_22 <= _zz_io_dataIn_0_payload_a_X_21;
    _zz_io_dataIn_0_payload_a_X_23 <= _zz_io_dataIn_0_payload_a_X_22;
    _zz_io_dataIn_0_payload_a_X_24 <= _zz_io_dataIn_0_payload_a_X_23;
    _zz_io_dataIn_0_payload_a_X_25 <= _zz_io_dataIn_0_payload_a_X_24;
    _zz_io_dataIn_0_payload_a_X_26 <= _zz_io_dataIn_0_payload_a_X_25;
    _zz_io_dataIn_0_payload_a_X_27 <= _zz_io_dataIn_0_payload_a_X_26;
    _zz_io_dataIn_0_payload_a_X_28 <= _zz_io_dataIn_0_payload_a_X_27;
    _zz_io_dataIn_0_payload_a_X_29 <= _zz_io_dataIn_0_payload_a_X_28;
    _zz_io_dataIn_0_payload_a_X_30 <= _zz_io_dataIn_0_payload_a_X_29;
    _zz_io_dataIn_0_payload_a_X_31 <= _zz_io_dataIn_0_payload_a_X_30;
    _zz_io_dataIn_0_payload_a_X_32 <= _zz_io_dataIn_0_payload_a_X_31;
    _zz_io_dataIn_0_payload_a_X_33 <= _zz_io_dataIn_0_payload_a_X_32;
    _zz_io_dataIn_0_payload_a_X_34 <= _zz_io_dataIn_0_payload_a_X_33;
    stage1_inputData_0_delay_1_X_1 <= stage1_inputData_0_X;
    stage1_inputData_0_delay_1_Y_1 <= stage1_inputData_0_Y;
    stage1_inputData_0_delay_1_Z_1 <= stage1_inputData_0_Z;
    stage1_inputData_0_delay_1_T_1 <= stage1_inputData_0_T;
    stage1_inputData_0_delay_2_X_1 <= stage1_inputData_0_delay_1_X_1;
    stage1_inputData_0_delay_2_Y_1 <= stage1_inputData_0_delay_1_Y_1;
    stage1_inputData_0_delay_2_Z_1 <= stage1_inputData_0_delay_1_Z_1;
    stage1_inputData_0_delay_2_T_1 <= stage1_inputData_0_delay_1_T_1;
    stage1_inputData_0_delay_3_X_1 <= stage1_inputData_0_delay_2_X_1;
    stage1_inputData_0_delay_3_Y_1 <= stage1_inputData_0_delay_2_Y_1;
    stage1_inputData_0_delay_3_Z_1 <= stage1_inputData_0_delay_2_Z_1;
    stage1_inputData_0_delay_3_T_1 <= stage1_inputData_0_delay_2_T_1;
    stage1_inputData_0_delay_4_X_1 <= stage1_inputData_0_delay_3_X_1;
    stage1_inputData_0_delay_4_Y_1 <= stage1_inputData_0_delay_3_Y_1;
    stage1_inputData_0_delay_4_Z_1 <= stage1_inputData_0_delay_3_Z_1;
    stage1_inputData_0_delay_4_T_1 <= stage1_inputData_0_delay_3_T_1;
    stage1_inputData_0_delay_5_X_1 <= stage1_inputData_0_delay_4_X_1;
    stage1_inputData_0_delay_5_Y_1 <= stage1_inputData_0_delay_4_Y_1;
    stage1_inputData_0_delay_5_Z_1 <= stage1_inputData_0_delay_4_Z_1;
    stage1_inputData_0_delay_5_T_1 <= stage1_inputData_0_delay_4_T_1;
    stage1_inputData_0_delay_6_X <= stage1_inputData_0_delay_5_X_1;
    stage1_inputData_0_delay_6_Y <= stage1_inputData_0_delay_5_Y_1;
    stage1_inputData_0_delay_6_Z <= stage1_inputData_0_delay_5_Z_1;
    stage1_inputData_0_delay_6_T <= stage1_inputData_0_delay_5_T_1;
    stage1_inputData_0_delay_7_X <= stage1_inputData_0_delay_6_X;
    stage1_inputData_0_delay_7_Y <= stage1_inputData_0_delay_6_Y;
    stage1_inputData_0_delay_7_Z <= stage1_inputData_0_delay_6_Z;
    stage1_inputData_0_delay_7_T <= stage1_inputData_0_delay_6_T;
    stage1_inputData_0_delay_8_X <= stage1_inputData_0_delay_7_X;
    stage1_inputData_0_delay_8_Y <= stage1_inputData_0_delay_7_Y;
    stage1_inputData_0_delay_8_Z <= stage1_inputData_0_delay_7_Z;
    stage1_inputData_0_delay_8_T <= stage1_inputData_0_delay_7_T;
    stage1_inputData_0_delay_9_X <= stage1_inputData_0_delay_8_X;
    stage1_inputData_0_delay_9_Y <= stage1_inputData_0_delay_8_Y;
    stage1_inputData_0_delay_9_Z <= stage1_inputData_0_delay_8_Z;
    stage1_inputData_0_delay_9_T <= stage1_inputData_0_delay_8_T;
    stage1_inputData_0_delay_10_X <= stage1_inputData_0_delay_9_X;
    stage1_inputData_0_delay_10_Y <= stage1_inputData_0_delay_9_Y;
    stage1_inputData_0_delay_10_Z <= stage1_inputData_0_delay_9_Z;
    stage1_inputData_0_delay_10_T <= stage1_inputData_0_delay_9_T;
    stage1_inputData_0_delay_11_X <= stage1_inputData_0_delay_10_X;
    stage1_inputData_0_delay_11_Y <= stage1_inputData_0_delay_10_Y;
    stage1_inputData_0_delay_11_Z <= stage1_inputData_0_delay_10_Z;
    stage1_inputData_0_delay_11_T <= stage1_inputData_0_delay_10_T;
    stage1_inputData_0_delay_12_X <= stage1_inputData_0_delay_11_X;
    stage1_inputData_0_delay_12_Y <= stage1_inputData_0_delay_11_Y;
    stage1_inputData_0_delay_12_Z <= stage1_inputData_0_delay_11_Z;
    stage1_inputData_0_delay_12_T <= stage1_inputData_0_delay_11_T;
    stage1_inputData_0_delay_13_X <= stage1_inputData_0_delay_12_X;
    stage1_inputData_0_delay_13_Y <= stage1_inputData_0_delay_12_Y;
    stage1_inputData_0_delay_13_Z <= stage1_inputData_0_delay_12_Z;
    stage1_inputData_0_delay_13_T <= stage1_inputData_0_delay_12_T;
    stage1_inputData_0_delay_14_X <= stage1_inputData_0_delay_13_X;
    stage1_inputData_0_delay_14_Y <= stage1_inputData_0_delay_13_Y;
    stage1_inputData_0_delay_14_Z <= stage1_inputData_0_delay_13_Z;
    stage1_inputData_0_delay_14_T <= stage1_inputData_0_delay_13_T;
    stage1_inputData_0_delay_15_X <= stage1_inputData_0_delay_14_X;
    stage1_inputData_0_delay_15_Y <= stage1_inputData_0_delay_14_Y;
    stage1_inputData_0_delay_15_Z <= stage1_inputData_0_delay_14_Z;
    stage1_inputData_0_delay_15_T <= stage1_inputData_0_delay_14_T;
    stage1_inputData_0_delay_16_X <= stage1_inputData_0_delay_15_X;
    stage1_inputData_0_delay_16_Y <= stage1_inputData_0_delay_15_Y;
    stage1_inputData_0_delay_16_Z <= stage1_inputData_0_delay_15_Z;
    stage1_inputData_0_delay_16_T <= stage1_inputData_0_delay_15_T;
    stage1_inputData_0_delay_17_X <= stage1_inputData_0_delay_16_X;
    stage1_inputData_0_delay_17_Y <= stage1_inputData_0_delay_16_Y;
    stage1_inputData_0_delay_17_Z <= stage1_inputData_0_delay_16_Z;
    stage1_inputData_0_delay_17_T <= stage1_inputData_0_delay_16_T;
    stage1_inputData_0_delay_18_X <= stage1_inputData_0_delay_17_X;
    stage1_inputData_0_delay_18_Y <= stage1_inputData_0_delay_17_Y;
    stage1_inputData_0_delay_18_Z <= stage1_inputData_0_delay_17_Z;
    stage1_inputData_0_delay_18_T <= stage1_inputData_0_delay_17_T;
    stage1_inputData_0_delay_19_X <= stage1_inputData_0_delay_18_X;
    stage1_inputData_0_delay_19_Y <= stage1_inputData_0_delay_18_Y;
    stage1_inputData_0_delay_19_Z <= stage1_inputData_0_delay_18_Z;
    stage1_inputData_0_delay_19_T <= stage1_inputData_0_delay_18_T;
    stage1_inputData_0_delay_20_X <= stage1_inputData_0_delay_19_X;
    stage1_inputData_0_delay_20_Y <= stage1_inputData_0_delay_19_Y;
    stage1_inputData_0_delay_20_Z <= stage1_inputData_0_delay_19_Z;
    stage1_inputData_0_delay_20_T <= stage1_inputData_0_delay_19_T;
    stage1_inputData_0_delay_21_X <= stage1_inputData_0_delay_20_X;
    stage1_inputData_0_delay_21_Y <= stage1_inputData_0_delay_20_Y;
    stage1_inputData_0_delay_21_Z <= stage1_inputData_0_delay_20_Z;
    stage1_inputData_0_delay_21_T <= stage1_inputData_0_delay_20_T;
    stage1_inputData_0_delay_22_X <= stage1_inputData_0_delay_21_X;
    stage1_inputData_0_delay_22_Y <= stage1_inputData_0_delay_21_Y;
    stage1_inputData_0_delay_22_Z <= stage1_inputData_0_delay_21_Z;
    stage1_inputData_0_delay_22_T <= stage1_inputData_0_delay_21_T;
    stage1_inputData_0_delay_23_X <= stage1_inputData_0_delay_22_X;
    stage1_inputData_0_delay_23_Y <= stage1_inputData_0_delay_22_Y;
    stage1_inputData_0_delay_23_Z <= stage1_inputData_0_delay_22_Z;
    stage1_inputData_0_delay_23_T <= stage1_inputData_0_delay_22_T;
    stage1_inputData_0_delay_24_X <= stage1_inputData_0_delay_23_X;
    stage1_inputData_0_delay_24_Y <= stage1_inputData_0_delay_23_Y;
    stage1_inputData_0_delay_24_Z <= stage1_inputData_0_delay_23_Z;
    stage1_inputData_0_delay_24_T <= stage1_inputData_0_delay_23_T;
    stage1_inputData_0_delay_25_X <= stage1_inputData_0_delay_24_X;
    stage1_inputData_0_delay_25_Y <= stage1_inputData_0_delay_24_Y;
    stage1_inputData_0_delay_25_Z <= stage1_inputData_0_delay_24_Z;
    stage1_inputData_0_delay_25_T <= stage1_inputData_0_delay_24_T;
    stage1_inputData_0_delay_26_X <= stage1_inputData_0_delay_25_X;
    stage1_inputData_0_delay_26_Y <= stage1_inputData_0_delay_25_Y;
    stage1_inputData_0_delay_26_Z <= stage1_inputData_0_delay_25_Z;
    stage1_inputData_0_delay_26_T <= stage1_inputData_0_delay_25_T;
    stage1_inputData_0_delay_27_X <= stage1_inputData_0_delay_26_X;
    stage1_inputData_0_delay_27_Y <= stage1_inputData_0_delay_26_Y;
    stage1_inputData_0_delay_27_Z <= stage1_inputData_0_delay_26_Z;
    stage1_inputData_0_delay_27_T <= stage1_inputData_0_delay_26_T;
    stage1_inputData_0_delay_28_X <= stage1_inputData_0_delay_27_X;
    stage1_inputData_0_delay_28_Y <= stage1_inputData_0_delay_27_Y;
    stage1_inputData_0_delay_28_Z <= stage1_inputData_0_delay_27_Z;
    stage1_inputData_0_delay_28_T <= stage1_inputData_0_delay_27_T;
    stage1_inputData_0_delay_29_X <= stage1_inputData_0_delay_28_X;
    stage1_inputData_0_delay_29_Y <= stage1_inputData_0_delay_28_Y;
    stage1_inputData_0_delay_29_Z <= stage1_inputData_0_delay_28_Z;
    stage1_inputData_0_delay_29_T <= stage1_inputData_0_delay_28_T;
    stage1_inputData_0_delay_30_X <= stage1_inputData_0_delay_29_X;
    stage1_inputData_0_delay_30_Y <= stage1_inputData_0_delay_29_Y;
    stage1_inputData_0_delay_30_Z <= stage1_inputData_0_delay_29_Z;
    stage1_inputData_0_delay_30_T <= stage1_inputData_0_delay_29_T;
    stage1_inputData_0_delay_31_X <= stage1_inputData_0_delay_30_X;
    stage1_inputData_0_delay_31_Y <= stage1_inputData_0_delay_30_Y;
    stage1_inputData_0_delay_31_Z <= stage1_inputData_0_delay_30_Z;
    stage1_inputData_0_delay_31_T <= stage1_inputData_0_delay_30_T;
    stage1_inputData_0_delay_32_X <= stage1_inputData_0_delay_31_X;
    stage1_inputData_0_delay_32_Y <= stage1_inputData_0_delay_31_Y;
    stage1_inputData_0_delay_32_Z <= stage1_inputData_0_delay_31_Z;
    stage1_inputData_0_delay_32_T <= stage1_inputData_0_delay_31_T;
    stage1_inputData_0_delay_33_X <= stage1_inputData_0_delay_32_X;
    stage1_inputData_0_delay_33_Y <= stage1_inputData_0_delay_32_Y;
    stage1_inputData_0_delay_33_Z <= stage1_inputData_0_delay_32_Z;
    stage1_inputData_0_delay_33_T <= stage1_inputData_0_delay_32_T;
    stage1_inputData_0_delay_34_X <= stage1_inputData_0_delay_33_X;
    stage1_inputData_0_delay_34_Y <= stage1_inputData_0_delay_33_Y;
    stage1_inputData_0_delay_34_Z <= stage1_inputData_0_delay_33_Z;
    stage1_inputData_0_delay_34_T <= stage1_inputData_0_delay_33_T;
    stage1_inputData_0_delay_35_X <= stage1_inputData_0_delay_34_X;
    stage1_inputData_0_delay_35_Y <= stage1_inputData_0_delay_34_Y;
    stage1_inputData_0_delay_35_Z <= stage1_inputData_0_delay_34_Z;
    stage1_inputData_0_delay_35_T <= stage1_inputData_0_delay_34_T;
    pAddPort_0_s_delay_1_X <= pAddPort_0_s_X;
    pAddPort_0_s_delay_1_Y <= pAddPort_0_s_Y;
    pAddPort_0_s_delay_1_Z <= pAddPort_0_s_Z;
    pAddPort_0_s_delay_1_T <= pAddPort_0_s_T;
    pAddPort_0_s_delay_2_X <= pAddPort_0_s_delay_1_X;
    pAddPort_0_s_delay_2_Y <= pAddPort_0_s_delay_1_Y;
    pAddPort_0_s_delay_2_Z <= pAddPort_0_s_delay_1_Z;
    pAddPort_0_s_delay_2_T <= pAddPort_0_s_delay_1_T;
    pAddPort_0_s_delay_3_X <= pAddPort_0_s_delay_2_X;
    pAddPort_0_s_delay_3_Y <= pAddPort_0_s_delay_2_Y;
    pAddPort_0_s_delay_3_Z <= pAddPort_0_s_delay_2_Z;
    pAddPort_0_s_delay_3_T <= pAddPort_0_s_delay_2_T;
    pAddPort_0_s_delay_4_X <= pAddPort_0_s_delay_3_X;
    pAddPort_0_s_delay_4_Y <= pAddPort_0_s_delay_3_Y;
    pAddPort_0_s_delay_4_Z <= pAddPort_0_s_delay_3_Z;
    pAddPort_0_s_delay_4_T <= pAddPort_0_s_delay_3_T;
    pAddPort_0_s_delay_5_X <= pAddPort_0_s_delay_4_X;
    pAddPort_0_s_delay_5_Y <= pAddPort_0_s_delay_4_Y;
    pAddPort_0_s_delay_5_Z <= pAddPort_0_s_delay_4_Z;
    pAddPort_0_s_delay_5_T <= pAddPort_0_s_delay_4_T;
    pAddPort_0_s_delay_6_X <= pAddPort_0_s_delay_5_X;
    pAddPort_0_s_delay_6_Y <= pAddPort_0_s_delay_5_Y;
    pAddPort_0_s_delay_6_Z <= pAddPort_0_s_delay_5_Z;
    pAddPort_0_s_delay_6_T <= pAddPort_0_s_delay_5_T;
    pAddPort_0_s_delay_7_X <= pAddPort_0_s_delay_6_X;
    pAddPort_0_s_delay_7_Y <= pAddPort_0_s_delay_6_Y;
    pAddPort_0_s_delay_7_Z <= pAddPort_0_s_delay_6_Z;
    pAddPort_0_s_delay_7_T <= pAddPort_0_s_delay_6_T;
    pAddPort_0_s_delay_8_X <= pAddPort_0_s_delay_7_X;
    pAddPort_0_s_delay_8_Y <= pAddPort_0_s_delay_7_Y;
    pAddPort_0_s_delay_8_Z <= pAddPort_0_s_delay_7_Z;
    pAddPort_0_s_delay_8_T <= pAddPort_0_s_delay_7_T;
    pAddPort_0_s_delay_9_X <= pAddPort_0_s_delay_8_X;
    pAddPort_0_s_delay_9_Y <= pAddPort_0_s_delay_8_Y;
    pAddPort_0_s_delay_9_Z <= pAddPort_0_s_delay_8_Z;
    pAddPort_0_s_delay_9_T <= pAddPort_0_s_delay_8_T;
    pAddPort_0_s_delay_10_X <= pAddPort_0_s_delay_9_X;
    pAddPort_0_s_delay_10_Y <= pAddPort_0_s_delay_9_Y;
    pAddPort_0_s_delay_10_Z <= pAddPort_0_s_delay_9_Z;
    pAddPort_0_s_delay_10_T <= pAddPort_0_s_delay_9_T;
    pAddPort_0_s_delay_11_X <= pAddPort_0_s_delay_10_X;
    pAddPort_0_s_delay_11_Y <= pAddPort_0_s_delay_10_Y;
    pAddPort_0_s_delay_11_Z <= pAddPort_0_s_delay_10_Z;
    pAddPort_0_s_delay_11_T <= pAddPort_0_s_delay_10_T;
    pAddPort_0_s_delay_12_X <= pAddPort_0_s_delay_11_X;
    pAddPort_0_s_delay_12_Y <= pAddPort_0_s_delay_11_Y;
    pAddPort_0_s_delay_12_Z <= pAddPort_0_s_delay_11_Z;
    pAddPort_0_s_delay_12_T <= pAddPort_0_s_delay_11_T;
    pAddPort_0_s_delay_13_X <= pAddPort_0_s_delay_12_X;
    pAddPort_0_s_delay_13_Y <= pAddPort_0_s_delay_12_Y;
    pAddPort_0_s_delay_13_Z <= pAddPort_0_s_delay_12_Z;
    pAddPort_0_s_delay_13_T <= pAddPort_0_s_delay_12_T;
    pAddPort_0_s_delay_14_X <= pAddPort_0_s_delay_13_X;
    pAddPort_0_s_delay_14_Y <= pAddPort_0_s_delay_13_Y;
    pAddPort_0_s_delay_14_Z <= pAddPort_0_s_delay_13_Z;
    pAddPort_0_s_delay_14_T <= pAddPort_0_s_delay_13_T;
    pAddPort_0_s_delay_15_X <= pAddPort_0_s_delay_14_X;
    pAddPort_0_s_delay_15_Y <= pAddPort_0_s_delay_14_Y;
    pAddPort_0_s_delay_15_Z <= pAddPort_0_s_delay_14_Z;
    pAddPort_0_s_delay_15_T <= pAddPort_0_s_delay_14_T;
    pAddPort_0_s_delay_16_X <= pAddPort_0_s_delay_15_X;
    pAddPort_0_s_delay_16_Y <= pAddPort_0_s_delay_15_Y;
    pAddPort_0_s_delay_16_Z <= pAddPort_0_s_delay_15_Z;
    pAddPort_0_s_delay_16_T <= pAddPort_0_s_delay_15_T;
    pAddPort_0_s_delay_17_X <= pAddPort_0_s_delay_16_X;
    pAddPort_0_s_delay_17_Y <= pAddPort_0_s_delay_16_Y;
    pAddPort_0_s_delay_17_Z <= pAddPort_0_s_delay_16_Z;
    pAddPort_0_s_delay_17_T <= pAddPort_0_s_delay_16_T;
    pAddPort_0_s_delay_18_X <= pAddPort_0_s_delay_17_X;
    pAddPort_0_s_delay_18_Y <= pAddPort_0_s_delay_17_Y;
    pAddPort_0_s_delay_18_Z <= pAddPort_0_s_delay_17_Z;
    pAddPort_0_s_delay_18_T <= pAddPort_0_s_delay_17_T;
    pAddPort_0_s_delay_19_X <= pAddPort_0_s_delay_18_X;
    pAddPort_0_s_delay_19_Y <= pAddPort_0_s_delay_18_Y;
    pAddPort_0_s_delay_19_Z <= pAddPort_0_s_delay_18_Z;
    pAddPort_0_s_delay_19_T <= pAddPort_0_s_delay_18_T;
    pAddPort_0_s_delay_20_X <= pAddPort_0_s_delay_19_X;
    pAddPort_0_s_delay_20_Y <= pAddPort_0_s_delay_19_Y;
    pAddPort_0_s_delay_20_Z <= pAddPort_0_s_delay_19_Z;
    pAddPort_0_s_delay_20_T <= pAddPort_0_s_delay_19_T;
    pAddPort_0_s_delay_21_X <= pAddPort_0_s_delay_20_X;
    pAddPort_0_s_delay_21_Y <= pAddPort_0_s_delay_20_Y;
    pAddPort_0_s_delay_21_Z <= pAddPort_0_s_delay_20_Z;
    pAddPort_0_s_delay_21_T <= pAddPort_0_s_delay_20_T;
    pAddPort_0_s_delay_22_X <= pAddPort_0_s_delay_21_X;
    pAddPort_0_s_delay_22_Y <= pAddPort_0_s_delay_21_Y;
    pAddPort_0_s_delay_22_Z <= pAddPort_0_s_delay_21_Z;
    pAddPort_0_s_delay_22_T <= pAddPort_0_s_delay_21_T;
    pAddPort_0_s_delay_23_X <= pAddPort_0_s_delay_22_X;
    pAddPort_0_s_delay_23_Y <= pAddPort_0_s_delay_22_Y;
    pAddPort_0_s_delay_23_Z <= pAddPort_0_s_delay_22_Z;
    pAddPort_0_s_delay_23_T <= pAddPort_0_s_delay_22_T;
    pAddPort_0_s_delay_24_X <= pAddPort_0_s_delay_23_X;
    pAddPort_0_s_delay_24_Y <= pAddPort_0_s_delay_23_Y;
    pAddPort_0_s_delay_24_Z <= pAddPort_0_s_delay_23_Z;
    pAddPort_0_s_delay_24_T <= pAddPort_0_s_delay_23_T;
    pAddPort_0_s_delay_25_X <= pAddPort_0_s_delay_24_X;
    pAddPort_0_s_delay_25_Y <= pAddPort_0_s_delay_24_Y;
    pAddPort_0_s_delay_25_Z <= pAddPort_0_s_delay_24_Z;
    pAddPort_0_s_delay_25_T <= pAddPort_0_s_delay_24_T;
    pAddPort_0_s_delay_26_X <= pAddPort_0_s_delay_25_X;
    pAddPort_0_s_delay_26_Y <= pAddPort_0_s_delay_25_Y;
    pAddPort_0_s_delay_26_Z <= pAddPort_0_s_delay_25_Z;
    pAddPort_0_s_delay_26_T <= pAddPort_0_s_delay_25_T;
    pAddPort_0_s_delay_27_X <= pAddPort_0_s_delay_26_X;
    pAddPort_0_s_delay_27_Y <= pAddPort_0_s_delay_26_Y;
    pAddPort_0_s_delay_27_Z <= pAddPort_0_s_delay_26_Z;
    pAddPort_0_s_delay_27_T <= pAddPort_0_s_delay_26_T;
    pAddPort_0_s_delay_28_X <= pAddPort_0_s_delay_27_X;
    pAddPort_0_s_delay_28_Y <= pAddPort_0_s_delay_27_Y;
    pAddPort_0_s_delay_28_Z <= pAddPort_0_s_delay_27_Z;
    pAddPort_0_s_delay_28_T <= pAddPort_0_s_delay_27_T;
    pAddPort_0_s_delay_29_X <= pAddPort_0_s_delay_28_X;
    pAddPort_0_s_delay_29_Y <= pAddPort_0_s_delay_28_Y;
    pAddPort_0_s_delay_29_Z <= pAddPort_0_s_delay_28_Z;
    pAddPort_0_s_delay_29_T <= pAddPort_0_s_delay_28_T;
    pAddPort_0_s_delay_30_X <= pAddPort_0_s_delay_29_X;
    pAddPort_0_s_delay_30_Y <= pAddPort_0_s_delay_29_Y;
    pAddPort_0_s_delay_30_Z <= pAddPort_0_s_delay_29_Z;
    pAddPort_0_s_delay_30_T <= pAddPort_0_s_delay_29_T;
    shiftRegs_addressOutFull_0_delay_1 <= shiftRegs_addressOutFull_0;
    shiftRegs_addressOutFull_0_delay_2 <= shiftRegs_addressOutFull_0_delay_1;
    shiftRegs_addressOutFull_0_delay_3 <= shiftRegs_addressOutFull_0_delay_2;
    shiftRegs_addressOutFull_0_delay_4 <= shiftRegs_addressOutFull_0_delay_3;
    shiftRegs_addressOutFull_0_delay_5 <= shiftRegs_addressOutFull_0_delay_4;
    shiftRegs_addressOutFull_0_delay_6 <= shiftRegs_addressOutFull_0_delay_5;
    shiftRegs_addressOutFull_0_delay_7 <= shiftRegs_addressOutFull_0_delay_6;
    shiftRegs_addressOutFull_0_delay_8 <= shiftRegs_addressOutFull_0_delay_7;
    shiftRegs_addressOutFull_0_delay_9 <= shiftRegs_addressOutFull_0_delay_8;
    shiftRegs_addressOutFull_0_delay_10 <= shiftRegs_addressOutFull_0_delay_9;
    shiftRegs_addressOutFull_0_delay_11 <= shiftRegs_addressOutFull_0_delay_10;
    shiftRegs_addressOutFull_0_delay_12 <= shiftRegs_addressOutFull_0_delay_11;
    shiftRegs_addressOutFull_0_delay_13 <= shiftRegs_addressOutFull_0_delay_12;
    shiftRegs_addressOutFull_0_delay_14 <= shiftRegs_addressOutFull_0_delay_13;
    shiftRegs_addressOutFull_0_delay_15 <= shiftRegs_addressOutFull_0_delay_14;
    shiftRegs_addressOutFull_0_delay_16 <= shiftRegs_addressOutFull_0_delay_15;
    shiftRegs_addressOutFull_0_delay_17 <= shiftRegs_addressOutFull_0_delay_16;
    shiftRegs_addressOutFull_0_delay_18 <= shiftRegs_addressOutFull_0_delay_17;
    shiftRegs_addressOutFull_0_delay_19 <= shiftRegs_addressOutFull_0_delay_18;
    shiftRegs_addressOutFull_0_delay_20 <= shiftRegs_addressOutFull_0_delay_19;
    shiftRegs_addressOutFull_0_delay_21 <= shiftRegs_addressOutFull_0_delay_20;
    shiftRegs_addressOutFull_0_delay_22 <= shiftRegs_addressOutFull_0_delay_21;
    shiftRegs_addressOutFull_0_delay_23 <= shiftRegs_addressOutFull_0_delay_22;
    shiftRegs_addressOutFull_0_delay_24 <= shiftRegs_addressOutFull_0_delay_23;
    shiftRegs_addressOutFull_0_delay_25 <= shiftRegs_addressOutFull_0_delay_24;
    shiftRegs_addressOutFull_0_delay_26 <= shiftRegs_addressOutFull_0_delay_25;
    shiftRegs_addressOutFull_0_delay_27 <= shiftRegs_addressOutFull_0_delay_26;
    shiftRegs_addressOutFull_0_delay_28 <= shiftRegs_addressOutFull_0_delay_27;
    shiftRegs_addressOutFull_0_delay_29 <= shiftRegs_addressOutFull_0_delay_28;
    shiftRegs_addressOutFull_0_delay_30 <= shiftRegs_addressOutFull_0_delay_29;
    stage1_inputData_0_delay_1_X_2 <= stage1_inputData_0_X;
    stage1_inputData_0_delay_1_Y_2 <= stage1_inputData_0_Y;
    stage1_inputData_0_delay_1_Z_2 <= stage1_inputData_0_Z;
    stage1_inputData_0_delay_1_T_2 <= stage1_inputData_0_T;
    stage1_inputData_0_delay_2_X_2 <= stage1_inputData_0_delay_1_X_2;
    stage1_inputData_0_delay_2_Y_2 <= stage1_inputData_0_delay_1_Y_2;
    stage1_inputData_0_delay_2_Z_2 <= stage1_inputData_0_delay_1_Z_2;
    stage1_inputData_0_delay_2_T_2 <= stage1_inputData_0_delay_1_T_2;
    stage1_inputData_0_delay_3_X_2 <= stage1_inputData_0_delay_2_X_2;
    stage1_inputData_0_delay_3_Y_2 <= stage1_inputData_0_delay_2_Y_2;
    stage1_inputData_0_delay_3_Z_2 <= stage1_inputData_0_delay_2_Z_2;
    stage1_inputData_0_delay_3_T_2 <= stage1_inputData_0_delay_2_T_2;
    stage1_inputData_0_delay_4_X_2 <= stage1_inputData_0_delay_3_X_2;
    stage1_inputData_0_delay_4_Y_2 <= stage1_inputData_0_delay_3_Y_2;
    stage1_inputData_0_delay_4_Z_2 <= stage1_inputData_0_delay_3_Z_2;
    stage1_inputData_0_delay_4_T_2 <= stage1_inputData_0_delay_3_T_2;
    stage1_inputData_0_delay_5_X_2 <= stage1_inputData_0_delay_4_X_2;
    stage1_inputData_0_delay_5_Y_2 <= stage1_inputData_0_delay_4_Y_2;
    stage1_inputData_0_delay_5_Z_2 <= stage1_inputData_0_delay_4_Z_2;
    stage1_inputData_0_delay_5_T_2 <= stage1_inputData_0_delay_4_T_2;
    stage1_inputData_0_delay_6_X_1 <= stage1_inputData_0_delay_5_X_2;
    stage1_inputData_0_delay_6_Y_1 <= stage1_inputData_0_delay_5_Y_2;
    stage1_inputData_0_delay_6_Z_1 <= stage1_inputData_0_delay_5_Z_2;
    stage1_inputData_0_delay_6_T_1 <= stage1_inputData_0_delay_5_T_2;
    stage1_inputData_0_delay_7_X_1 <= stage1_inputData_0_delay_6_X_1;
    stage1_inputData_0_delay_7_Y_1 <= stage1_inputData_0_delay_6_Y_1;
    stage1_inputData_0_delay_7_Z_1 <= stage1_inputData_0_delay_6_Z_1;
    stage1_inputData_0_delay_7_T_1 <= stage1_inputData_0_delay_6_T_1;
    stage1_inputData_0_delay_8_X_1 <= stage1_inputData_0_delay_7_X_1;
    stage1_inputData_0_delay_8_Y_1 <= stage1_inputData_0_delay_7_Y_1;
    stage1_inputData_0_delay_8_Z_1 <= stage1_inputData_0_delay_7_Z_1;
    stage1_inputData_0_delay_8_T_1 <= stage1_inputData_0_delay_7_T_1;
    stage1_inputData_0_delay_9_X_1 <= stage1_inputData_0_delay_8_X_1;
    stage1_inputData_0_delay_9_Y_1 <= stage1_inputData_0_delay_8_Y_1;
    stage1_inputData_0_delay_9_Z_1 <= stage1_inputData_0_delay_8_Z_1;
    stage1_inputData_0_delay_9_T_1 <= stage1_inputData_0_delay_8_T_1;
    stage1_inputData_0_delay_10_X_1 <= stage1_inputData_0_delay_9_X_1;
    stage1_inputData_0_delay_10_Y_1 <= stage1_inputData_0_delay_9_Y_1;
    stage1_inputData_0_delay_10_Z_1 <= stage1_inputData_0_delay_9_Z_1;
    stage1_inputData_0_delay_10_T_1 <= stage1_inputData_0_delay_9_T_1;
    stage1_inputData_0_delay_11_X_1 <= stage1_inputData_0_delay_10_X_1;
    stage1_inputData_0_delay_11_Y_1 <= stage1_inputData_0_delay_10_Y_1;
    stage1_inputData_0_delay_11_Z_1 <= stage1_inputData_0_delay_10_Z_1;
    stage1_inputData_0_delay_11_T_1 <= stage1_inputData_0_delay_10_T_1;
    stage1_inputData_0_delay_12_X_1 <= stage1_inputData_0_delay_11_X_1;
    stage1_inputData_0_delay_12_Y_1 <= stage1_inputData_0_delay_11_Y_1;
    stage1_inputData_0_delay_12_Z_1 <= stage1_inputData_0_delay_11_Z_1;
    stage1_inputData_0_delay_12_T_1 <= stage1_inputData_0_delay_11_T_1;
    stage1_inputData_0_delay_13_X_1 <= stage1_inputData_0_delay_12_X_1;
    stage1_inputData_0_delay_13_Y_1 <= stage1_inputData_0_delay_12_Y_1;
    stage1_inputData_0_delay_13_Z_1 <= stage1_inputData_0_delay_12_Z_1;
    stage1_inputData_0_delay_13_T_1 <= stage1_inputData_0_delay_12_T_1;
    stage1_inputData_0_delay_14_X_1 <= stage1_inputData_0_delay_13_X_1;
    stage1_inputData_0_delay_14_Y_1 <= stage1_inputData_0_delay_13_Y_1;
    stage1_inputData_0_delay_14_Z_1 <= stage1_inputData_0_delay_13_Z_1;
    stage1_inputData_0_delay_14_T_1 <= stage1_inputData_0_delay_13_T_1;
    stage1_inputData_0_delay_15_X_1 <= stage1_inputData_0_delay_14_X_1;
    stage1_inputData_0_delay_15_Y_1 <= stage1_inputData_0_delay_14_Y_1;
    stage1_inputData_0_delay_15_Z_1 <= stage1_inputData_0_delay_14_Z_1;
    stage1_inputData_0_delay_15_T_1 <= stage1_inputData_0_delay_14_T_1;
    stage1_inputData_0_delay_16_X_1 <= stage1_inputData_0_delay_15_X_1;
    stage1_inputData_0_delay_16_Y_1 <= stage1_inputData_0_delay_15_Y_1;
    stage1_inputData_0_delay_16_Z_1 <= stage1_inputData_0_delay_15_Z_1;
    stage1_inputData_0_delay_16_T_1 <= stage1_inputData_0_delay_15_T_1;
    stage1_inputData_0_delay_17_X_1 <= stage1_inputData_0_delay_16_X_1;
    stage1_inputData_0_delay_17_Y_1 <= stage1_inputData_0_delay_16_Y_1;
    stage1_inputData_0_delay_17_Z_1 <= stage1_inputData_0_delay_16_Z_1;
    stage1_inputData_0_delay_17_T_1 <= stage1_inputData_0_delay_16_T_1;
    stage1_inputData_0_delay_18_X_1 <= stage1_inputData_0_delay_17_X_1;
    stage1_inputData_0_delay_18_Y_1 <= stage1_inputData_0_delay_17_Y_1;
    stage1_inputData_0_delay_18_Z_1 <= stage1_inputData_0_delay_17_Z_1;
    stage1_inputData_0_delay_18_T_1 <= stage1_inputData_0_delay_17_T_1;
    stage1_inputData_0_delay_19_X_1 <= stage1_inputData_0_delay_18_X_1;
    stage1_inputData_0_delay_19_Y_1 <= stage1_inputData_0_delay_18_Y_1;
    stage1_inputData_0_delay_19_Z_1 <= stage1_inputData_0_delay_18_Z_1;
    stage1_inputData_0_delay_19_T_1 <= stage1_inputData_0_delay_18_T_1;
    stage1_inputData_0_delay_20_X_1 <= stage1_inputData_0_delay_19_X_1;
    stage1_inputData_0_delay_20_Y_1 <= stage1_inputData_0_delay_19_Y_1;
    stage1_inputData_0_delay_20_Z_1 <= stage1_inputData_0_delay_19_Z_1;
    stage1_inputData_0_delay_20_T_1 <= stage1_inputData_0_delay_19_T_1;
    stage1_inputData_0_delay_21_X_1 <= stage1_inputData_0_delay_20_X_1;
    stage1_inputData_0_delay_21_Y_1 <= stage1_inputData_0_delay_20_Y_1;
    stage1_inputData_0_delay_21_Z_1 <= stage1_inputData_0_delay_20_Z_1;
    stage1_inputData_0_delay_21_T_1 <= stage1_inputData_0_delay_20_T_1;
    stage1_inputData_0_delay_22_X_1 <= stage1_inputData_0_delay_21_X_1;
    stage1_inputData_0_delay_22_Y_1 <= stage1_inputData_0_delay_21_Y_1;
    stage1_inputData_0_delay_22_Z_1 <= stage1_inputData_0_delay_21_Z_1;
    stage1_inputData_0_delay_22_T_1 <= stage1_inputData_0_delay_21_T_1;
    stage1_inputData_0_delay_23_X_1 <= stage1_inputData_0_delay_22_X_1;
    stage1_inputData_0_delay_23_Y_1 <= stage1_inputData_0_delay_22_Y_1;
    stage1_inputData_0_delay_23_Z_1 <= stage1_inputData_0_delay_22_Z_1;
    stage1_inputData_0_delay_23_T_1 <= stage1_inputData_0_delay_22_T_1;
    stage1_inputData_0_delay_24_X_1 <= stage1_inputData_0_delay_23_X_1;
    stage1_inputData_0_delay_24_Y_1 <= stage1_inputData_0_delay_23_Y_1;
    stage1_inputData_0_delay_24_Z_1 <= stage1_inputData_0_delay_23_Z_1;
    stage1_inputData_0_delay_24_T_1 <= stage1_inputData_0_delay_23_T_1;
    stage1_inputData_0_delay_25_X_1 <= stage1_inputData_0_delay_24_X_1;
    stage1_inputData_0_delay_25_Y_1 <= stage1_inputData_0_delay_24_Y_1;
    stage1_inputData_0_delay_25_Z_1 <= stage1_inputData_0_delay_24_Z_1;
    stage1_inputData_0_delay_25_T_1 <= stage1_inputData_0_delay_24_T_1;
    stage1_inputData_0_delay_26_X_1 <= stage1_inputData_0_delay_25_X_1;
    stage1_inputData_0_delay_26_Y_1 <= stage1_inputData_0_delay_25_Y_1;
    stage1_inputData_0_delay_26_Z_1 <= stage1_inputData_0_delay_25_Z_1;
    stage1_inputData_0_delay_26_T_1 <= stage1_inputData_0_delay_25_T_1;
    stage1_inputData_0_delay_27_X_1 <= stage1_inputData_0_delay_26_X_1;
    stage1_inputData_0_delay_27_Y_1 <= stage1_inputData_0_delay_26_Y_1;
    stage1_inputData_0_delay_27_Z_1 <= stage1_inputData_0_delay_26_Z_1;
    stage1_inputData_0_delay_27_T_1 <= stage1_inputData_0_delay_26_T_1;
    stage1_inputData_0_delay_28_X_1 <= stage1_inputData_0_delay_27_X_1;
    stage1_inputData_0_delay_28_Y_1 <= stage1_inputData_0_delay_27_Y_1;
    stage1_inputData_0_delay_28_Z_1 <= stage1_inputData_0_delay_27_Z_1;
    stage1_inputData_0_delay_28_T_1 <= stage1_inputData_0_delay_27_T_1;
    stage1_inputData_0_delay_29_X_1 <= stage1_inputData_0_delay_28_X_1;
    stage1_inputData_0_delay_29_Y_1 <= stage1_inputData_0_delay_28_Y_1;
    stage1_inputData_0_delay_29_Z_1 <= stage1_inputData_0_delay_28_Z_1;
    stage1_inputData_0_delay_29_T_1 <= stage1_inputData_0_delay_28_T_1;
    stage1_inputData_0_delay_30_X_1 <= stage1_inputData_0_delay_29_X_1;
    stage1_inputData_0_delay_30_Y_1 <= stage1_inputData_0_delay_29_Y_1;
    stage1_inputData_0_delay_30_Z_1 <= stage1_inputData_0_delay_29_Z_1;
    stage1_inputData_0_delay_30_T_1 <= stage1_inputData_0_delay_29_T_1;
    stage1_inputData_0_delay_31_X_1 <= stage1_inputData_0_delay_30_X_1;
    stage1_inputData_0_delay_31_Y_1 <= stage1_inputData_0_delay_30_Y_1;
    stage1_inputData_0_delay_31_Z_1 <= stage1_inputData_0_delay_30_Z_1;
    stage1_inputData_0_delay_31_T_1 <= stage1_inputData_0_delay_30_T_1;
    stage1_inputData_0_delay_32_X_1 <= stage1_inputData_0_delay_31_X_1;
    stage1_inputData_0_delay_32_Y_1 <= stage1_inputData_0_delay_31_Y_1;
    stage1_inputData_0_delay_32_Z_1 <= stage1_inputData_0_delay_31_Z_1;
    stage1_inputData_0_delay_32_T_1 <= stage1_inputData_0_delay_31_T_1;
    stage1_inputData_0_delay_33_X_1 <= stage1_inputData_0_delay_32_X_1;
    stage1_inputData_0_delay_33_Y_1 <= stage1_inputData_0_delay_32_Y_1;
    stage1_inputData_0_delay_33_Z_1 <= stage1_inputData_0_delay_32_Z_1;
    stage1_inputData_0_delay_33_T_1 <= stage1_inputData_0_delay_32_T_1;
    stage1_inputData_0_delay_34_X_1 <= stage1_inputData_0_delay_33_X_1;
    stage1_inputData_0_delay_34_Y_1 <= stage1_inputData_0_delay_33_Y_1;
    stage1_inputData_0_delay_34_Z_1 <= stage1_inputData_0_delay_33_Z_1;
    stage1_inputData_0_delay_34_T_1 <= stage1_inputData_0_delay_33_T_1;
    stage1_inputData_0_delay_35_X_1 <= stage1_inputData_0_delay_34_X_1;
    stage1_inputData_0_delay_35_Y_1 <= stage1_inputData_0_delay_34_Y_1;
    stage1_inputData_0_delay_35_Z_1 <= stage1_inputData_0_delay_34_Z_1;
    stage1_inputData_0_delay_35_T_1 <= stage1_inputData_0_delay_34_T_1;
    stage1_inputAddress_0_delay_1_1 <= stage1_inputAddress_0;
    stage1_inputAddress_0_delay_2_1 <= stage1_inputAddress_0_delay_1_1;
    stage1_inputAddress_0_delay_3_1 <= stage1_inputAddress_0_delay_2_1;
    stage1_inputAddress_0_delay_4_1 <= stage1_inputAddress_0_delay_3_1;
    stage1_inputAddress_0_delay_5_1 <= stage1_inputAddress_0_delay_4_1;
    stage1_inputAddress_0_delay_6 <= stage1_inputAddress_0_delay_5_1;
    stage1_inputAddress_0_delay_7 <= stage1_inputAddress_0_delay_6;
    stage1_inputAddress_0_delay_8 <= stage1_inputAddress_0_delay_7;
    stage1_inputAddress_0_delay_9 <= stage1_inputAddress_0_delay_8;
    stage1_inputAddress_0_delay_10 <= stage1_inputAddress_0_delay_9;
    stage1_inputAddress_0_delay_11 <= stage1_inputAddress_0_delay_10;
    stage1_inputAddress_0_delay_12 <= stage1_inputAddress_0_delay_11;
    stage1_inputAddress_0_delay_13 <= stage1_inputAddress_0_delay_12;
    stage1_inputAddress_0_delay_14 <= stage1_inputAddress_0_delay_13;
    stage1_inputAddress_0_delay_15 <= stage1_inputAddress_0_delay_14;
    stage1_inputAddress_0_delay_16 <= stage1_inputAddress_0_delay_15;
    stage1_inputAddress_0_delay_17 <= stage1_inputAddress_0_delay_16;
    stage1_inputAddress_0_delay_18 <= stage1_inputAddress_0_delay_17;
    stage1_inputAddress_0_delay_19 <= stage1_inputAddress_0_delay_18;
    stage1_inputAddress_0_delay_20 <= stage1_inputAddress_0_delay_19;
    stage1_inputAddress_0_delay_21 <= stage1_inputAddress_0_delay_20;
    stage1_inputAddress_0_delay_22 <= stage1_inputAddress_0_delay_21;
    stage1_inputAddress_0_delay_23 <= stage1_inputAddress_0_delay_22;
    stage1_inputAddress_0_delay_24 <= stage1_inputAddress_0_delay_23;
    stage1_inputAddress_0_delay_25 <= stage1_inputAddress_0_delay_24;
    stage1_inputAddress_0_delay_26 <= stage1_inputAddress_0_delay_25;
    stage1_inputAddress_0_delay_27 <= stage1_inputAddress_0_delay_26;
    stage1_inputAddress_0_delay_28 <= stage1_inputAddress_0_delay_27;
    stage1_inputAddress_0_delay_29 <= stage1_inputAddress_0_delay_28;
    stage1_inputAddress_0_delay_30 <= stage1_inputAddress_0_delay_29;
    stage1_inputAddress_0_delay_31 <= stage1_inputAddress_0_delay_30;
    stage1_inputAddress_0_delay_32 <= stage1_inputAddress_0_delay_31;
    stage1_inputAddress_0_delay_33 <= stage1_inputAddress_0_delay_32;
    stage1_inputAddress_0_delay_34 <= stage1_inputAddress_0_delay_33;
    stage1_inputAddress_0_delay_35 <= stage1_inputAddress_0_delay_34;
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      _zz_io_dataIn_0_valid_5 <= 1'b0;
      _zz_io_dataIn_0_valid_6 <= 1'b0;
      _zz_io_dataIn_0_valid_7 <= 1'b0;
      _zz_io_dataIn_0_valid_8 <= 1'b0;
      _zz_io_dataIn_0_valid_9 <= 1'b0;
      _zz_io_dataIn_0_valid_10 <= 1'b0;
      _zz_io_dataIn_0_valid_11 <= 1'b0;
      _zz_io_dataIn_0_valid_12 <= 1'b0;
      _zz_io_dataIn_0_valid_13 <= 1'b0;
      _zz_io_dataIn_0_valid_14 <= 1'b0;
      _zz_io_dataIn_0_valid_15 <= 1'b0;
      _zz_io_dataIn_0_valid_16 <= 1'b0;
      _zz_io_dataIn_0_valid_17 <= 1'b0;
      _zz_io_dataIn_0_valid_18 <= 1'b0;
      _zz_io_dataIn_0_valid_19 <= 1'b0;
      _zz_io_dataIn_0_valid_20 <= 1'b0;
      _zz_io_dataIn_0_valid_21 <= 1'b0;
      _zz_io_dataIn_0_valid_22 <= 1'b0;
      _zz_io_dataIn_0_valid_23 <= 1'b0;
      _zz_io_dataIn_0_valid_24 <= 1'b0;
      _zz_io_dataIn_0_valid_25 <= 1'b0;
      _zz_io_dataIn_0_valid_26 <= 1'b0;
      _zz_io_dataIn_0_valid_27 <= 1'b0;
      _zz_io_dataIn_0_valid_28 <= 1'b0;
      _zz_io_dataIn_0_valid_29 <= 1'b0;
      _zz_io_dataIn_0_valid_30 <= 1'b0;
      _zz_io_dataIn_0_valid_31 <= 1'b0;
      _zz_io_dataIn_0_valid_32 <= 1'b0;
      _zz_io_dataIn_0_valid_33 <= 1'b0;
      _zz_io_dataIn_0_valid_34 <= 1'b0;
      _zz_io_dataIn_1_valid <= 1'b0;
      _zz_io_dataIn_1_valid_1 <= 1'b0;
      _zz_io_dataIn_1_valid_2 <= 1'b0;
      _zz_io_dataIn_1_valid_3 <= 1'b0;
      _zz_io_dataIn_1_valid_4 <= 1'b0;
      _zz_io_dataIn_1_valid_5 <= 1'b0;
      _zz_io_dataIn_1_valid_6 <= 1'b0;
      _zz_io_dataIn_1_valid_7 <= 1'b0;
      _zz_io_dataIn_1_valid_8 <= 1'b0;
      _zz_io_dataIn_1_valid_9 <= 1'b0;
      _zz_io_dataIn_1_valid_10 <= 1'b0;
      _zz_io_dataIn_1_valid_11 <= 1'b0;
      _zz_io_dataIn_1_valid_12 <= 1'b0;
      _zz_io_dataIn_1_valid_13 <= 1'b0;
      _zz_io_dataIn_1_valid_14 <= 1'b0;
      _zz_io_dataIn_1_valid_15 <= 1'b0;
      _zz_io_dataIn_1_valid_16 <= 1'b0;
      _zz_io_dataIn_1_valid_17 <= 1'b0;
      _zz_io_dataIn_1_valid_18 <= 1'b0;
      _zz_io_dataIn_1_valid_19 <= 1'b0;
      _zz_io_dataIn_1_valid_20 <= 1'b0;
      _zz_io_dataIn_1_valid_21 <= 1'b0;
      _zz_io_dataIn_1_valid_22 <= 1'b0;
      _zz_io_dataIn_1_valid_23 <= 1'b0;
      _zz_io_dataIn_1_valid_24 <= 1'b0;
      _zz_io_dataIn_1_valid_25 <= 1'b0;
      _zz_io_dataIn_1_valid_26 <= 1'b0;
      _zz_io_dataIn_1_valid_27 <= 1'b0;
      _zz_io_dataIn_1_valid_28 <= 1'b0;
      _zz_io_dataIn_1_valid_29 <= 1'b0;
      _zz_io_dataIn_1_valid_30 <= 1'b0;
      _zz_io_dataIn_1_valid_31 <= 1'b0;
      _zz_io_dataIn_1_valid_32 <= 1'b0;
      _zz_io_dataIn_1_valid_33 <= 1'b0;
      _zz_io_dataIn_1_valid_34 <= 1'b0;
    end else begin
      _zz_io_dataIn_0_valid_5 <= ((stateRam_0_io_state_0 || _zz_io_dataIn_0_valid_4) && shiftRegs_validOutFull_0);
      _zz_io_dataIn_0_valid_6 <= _zz_io_dataIn_0_valid_5;
      _zz_io_dataIn_0_valid_7 <= _zz_io_dataIn_0_valid_6;
      _zz_io_dataIn_0_valid_8 <= _zz_io_dataIn_0_valid_7;
      _zz_io_dataIn_0_valid_9 <= _zz_io_dataIn_0_valid_8;
      _zz_io_dataIn_0_valid_10 <= _zz_io_dataIn_0_valid_9;
      _zz_io_dataIn_0_valid_11 <= _zz_io_dataIn_0_valid_10;
      _zz_io_dataIn_0_valid_12 <= _zz_io_dataIn_0_valid_11;
      _zz_io_dataIn_0_valid_13 <= _zz_io_dataIn_0_valid_12;
      _zz_io_dataIn_0_valid_14 <= _zz_io_dataIn_0_valid_13;
      _zz_io_dataIn_0_valid_15 <= _zz_io_dataIn_0_valid_14;
      _zz_io_dataIn_0_valid_16 <= _zz_io_dataIn_0_valid_15;
      _zz_io_dataIn_0_valid_17 <= _zz_io_dataIn_0_valid_16;
      _zz_io_dataIn_0_valid_18 <= _zz_io_dataIn_0_valid_17;
      _zz_io_dataIn_0_valid_19 <= _zz_io_dataIn_0_valid_18;
      _zz_io_dataIn_0_valid_20 <= _zz_io_dataIn_0_valid_19;
      _zz_io_dataIn_0_valid_21 <= _zz_io_dataIn_0_valid_20;
      _zz_io_dataIn_0_valid_22 <= _zz_io_dataIn_0_valid_21;
      _zz_io_dataIn_0_valid_23 <= _zz_io_dataIn_0_valid_22;
      _zz_io_dataIn_0_valid_24 <= _zz_io_dataIn_0_valid_23;
      _zz_io_dataIn_0_valid_25 <= _zz_io_dataIn_0_valid_24;
      _zz_io_dataIn_0_valid_26 <= _zz_io_dataIn_0_valid_25;
      _zz_io_dataIn_0_valid_27 <= _zz_io_dataIn_0_valid_26;
      _zz_io_dataIn_0_valid_28 <= _zz_io_dataIn_0_valid_27;
      _zz_io_dataIn_0_valid_29 <= _zz_io_dataIn_0_valid_28;
      _zz_io_dataIn_0_valid_30 <= _zz_io_dataIn_0_valid_29;
      _zz_io_dataIn_0_valid_31 <= _zz_io_dataIn_0_valid_30;
      _zz_io_dataIn_0_valid_32 <= _zz_io_dataIn_0_valid_31;
      _zz_io_dataIn_0_valid_33 <= _zz_io_dataIn_0_valid_32;
      _zz_io_dataIn_0_valid_34 <= _zz_io_dataIn_0_valid_33;
      _zz_io_dataIn_1_valid <= (stage1_inputValid_0 && (! (shiftRegs_validOut_0 && (stage1_inputAddress_0 == shiftRegs_addressOut_0))));
      _zz_io_dataIn_1_valid_1 <= _zz_io_dataIn_1_valid;
      _zz_io_dataIn_1_valid_2 <= _zz_io_dataIn_1_valid_1;
      _zz_io_dataIn_1_valid_3 <= _zz_io_dataIn_1_valid_2;
      _zz_io_dataIn_1_valid_4 <= _zz_io_dataIn_1_valid_3;
      _zz_io_dataIn_1_valid_5 <= (stateRam_0_io_state_1 && _zz_io_dataIn_1_valid_4);
      _zz_io_dataIn_1_valid_6 <= _zz_io_dataIn_1_valid_5;
      _zz_io_dataIn_1_valid_7 <= _zz_io_dataIn_1_valid_6;
      _zz_io_dataIn_1_valid_8 <= _zz_io_dataIn_1_valid_7;
      _zz_io_dataIn_1_valid_9 <= _zz_io_dataIn_1_valid_8;
      _zz_io_dataIn_1_valid_10 <= _zz_io_dataIn_1_valid_9;
      _zz_io_dataIn_1_valid_11 <= _zz_io_dataIn_1_valid_10;
      _zz_io_dataIn_1_valid_12 <= _zz_io_dataIn_1_valid_11;
      _zz_io_dataIn_1_valid_13 <= _zz_io_dataIn_1_valid_12;
      _zz_io_dataIn_1_valid_14 <= _zz_io_dataIn_1_valid_13;
      _zz_io_dataIn_1_valid_15 <= _zz_io_dataIn_1_valid_14;
      _zz_io_dataIn_1_valid_16 <= _zz_io_dataIn_1_valid_15;
      _zz_io_dataIn_1_valid_17 <= _zz_io_dataIn_1_valid_16;
      _zz_io_dataIn_1_valid_18 <= _zz_io_dataIn_1_valid_17;
      _zz_io_dataIn_1_valid_19 <= _zz_io_dataIn_1_valid_18;
      _zz_io_dataIn_1_valid_20 <= _zz_io_dataIn_1_valid_19;
      _zz_io_dataIn_1_valid_21 <= _zz_io_dataIn_1_valid_20;
      _zz_io_dataIn_1_valid_22 <= _zz_io_dataIn_1_valid_21;
      _zz_io_dataIn_1_valid_23 <= _zz_io_dataIn_1_valid_22;
      _zz_io_dataIn_1_valid_24 <= _zz_io_dataIn_1_valid_23;
      _zz_io_dataIn_1_valid_25 <= _zz_io_dataIn_1_valid_24;
      _zz_io_dataIn_1_valid_26 <= _zz_io_dataIn_1_valid_25;
      _zz_io_dataIn_1_valid_27 <= _zz_io_dataIn_1_valid_26;
      _zz_io_dataIn_1_valid_28 <= _zz_io_dataIn_1_valid_27;
      _zz_io_dataIn_1_valid_29 <= _zz_io_dataIn_1_valid_28;
      _zz_io_dataIn_1_valid_30 <= _zz_io_dataIn_1_valid_29;
      _zz_io_dataIn_1_valid_31 <= _zz_io_dataIn_1_valid_30;
      _zz_io_dataIn_1_valid_32 <= _zz_io_dataIn_1_valid_31;
      _zz_io_dataIn_1_valid_33 <= _zz_io_dataIn_1_valid_32;
      _zz_io_dataIn_1_valid_34 <= _zz_io_dataIn_1_valid_33;
    end
  end

  always @(posedge clk) begin
    _zz_io_state_1 <= (stage2_wCnt_value == 12'hfff);
    _zz_io_state_1_1 <= _zz_io_state_1;
    _zz_io_state_1_2 <= _zz_io_state_1_1;
    _zz_io_state_1_3 <= _zz_io_state_1_2;
    _zz_io_state_1_4 <= _zz_io_state_1_3;
    _zz_io_state_1_5 <= (! stage2_calCnt_value[1]);
    _zz_io_state_1_6 <= _zz_io_state_1_5;
    _zz_io_state_1_7 <= _zz_io_state_1_6;
    _zz_io_state_1_8 <= _zz_io_state_1_7;
    _zz_io_state_1_9 <= _zz_io_state_1_8;
    _zz_io_state_1_10 <= (|stage2_calCnt_value);
    _zz_io_state_1_11 <= _zz_io_state_1_10;
    _zz_io_state_1_12 <= _zz_io_state_1_11;
    _zz_io_state_1_13 <= _zz_io_state_1_12;
    _zz_io_state_1_14 <= _zz_io_state_1_13;
    _zz_io_state_1_15 <= (_zz_io_state_1_4 ? (_zz_io_state_1_9 && stateRam_0_io_state_0) : (_zz_io_state_1_14 || stateRam_0_io_state_0));
    _zz_io_state_1_16 <= _zz_io_state_1_15;
    _zz_io_state_1_17 <= _zz_io_state_1_16;
    _zz_io_state_1_18 <= _zz_io_state_1_17;
    _zz_io_state_1_19 <= _zz_io_state_1_18;
    _zz_io_state_1_20 <= _zz_io_state_1_19;
    _zz_io_state_1_21 <= _zz_io_state_1_20;
    _zz_io_state_1_22 <= _zz_io_state_1_21;
    _zz_io_state_1_23 <= _zz_io_state_1_22;
    _zz_io_state_1_24 <= _zz_io_state_1_23;
    _zz_io_state_1_25 <= _zz_io_state_1_24;
    _zz_io_state_1_26 <= _zz_io_state_1_25;
    _zz_io_state_1_27 <= _zz_io_state_1_26;
    _zz_io_state_1_28 <= _zz_io_state_1_27;
    _zz_io_state_1_29 <= _zz_io_state_1_28;
    _zz_io_state_1_30 <= _zz_io_state_1_29;
    _zz_io_state_1_31 <= _zz_io_state_1_30;
    _zz_io_state_1_32 <= _zz_io_state_1_31;
    _zz_io_state_1_33 <= _zz_io_state_1_32;
    _zz_io_state_1_34 <= _zz_io_state_1_33;
    _zz_io_state_1_35 <= _zz_io_state_1_34;
    _zz_io_state_1_36 <= _zz_io_state_1_35;
    _zz_io_state_1_37 <= _zz_io_state_1_36;
    _zz_io_state_1_38 <= _zz_io_state_1_37;
    pippenger_1_dataRam_0_io_rData_1_regNext_X <= dataRam_0_io_rData_1_X;
    pippenger_1_dataRam_0_io_rData_1_regNext_Y <= dataRam_0_io_rData_1_Y;
    pippenger_1_dataRam_0_io_rData_1_regNext_Z <= dataRam_0_io_rData_1_Z;
    pippenger_1_dataRam_0_io_rData_1_regNext_T <= dataRam_0_io_rData_1_T;
    _zz_io_dataIn_1_payload_address <= {stage2_GCnt_value,_zz__zz_io_dataIn_1_payload_address};
    _zz_io_dataIn_1_payload_address_1 <= _zz_io_dataIn_1_payload_address;
    _zz_io_dataIn_1_payload_address_2 <= _zz_io_dataIn_1_payload_address_1;
    _zz_io_dataIn_1_payload_address_3 <= _zz_io_dataIn_1_payload_address_2;
    _zz_io_dataIn_1_payload_address_4 <= _zz_io_dataIn_1_payload_address_3;
    _zz_io_dataIn_1_payload_address_5 <= _zz_io_dataIn_1_payload_address_4;
    _zz_io_dataIn_1_payload_address_6 <= _zz_io_dataIn_1_payload_address_5;
    _zz_io_dataIn_1_payload_address_7 <= _zz_io_dataIn_1_payload_address_6;
    _zz_io_dataIn_1_payload_address_8 <= _zz_io_dataIn_1_payload_address_7;
    _zz_io_dataIn_1_payload_address_9 <= _zz_io_dataIn_1_payload_address_8;
    _zz_io_dataIn_1_payload_address_10 <= _zz_io_dataIn_1_payload_address_9;
    _zz_io_dataIn_1_payload_address_11 <= _zz_io_dataIn_1_payload_address_10;
    _zz_io_dataIn_1_payload_address_12 <= _zz_io_dataIn_1_payload_address_11;
    _zz_io_dataIn_1_payload_address_13 <= _zz_io_dataIn_1_payload_address_12;
    _zz_io_dataIn_1_payload_address_14 <= _zz_io_dataIn_1_payload_address_13;
    _zz_io_dataIn_1_payload_address_15 <= _zz_io_dataIn_1_payload_address_14;
    _zz_io_dataIn_1_payload_address_16 <= _zz_io_dataIn_1_payload_address_15;
    _zz_io_dataIn_1_payload_address_17 <= _zz_io_dataIn_1_payload_address_16;
    _zz_io_dataIn_1_payload_address_18 <= _zz_io_dataIn_1_payload_address_17;
    _zz_io_dataIn_1_payload_address_19 <= _zz_io_dataIn_1_payload_address_18;
    _zz_io_dataIn_1_payload_address_20 <= _zz_io_dataIn_1_payload_address_19;
    _zz_io_dataIn_1_payload_address_21 <= _zz_io_dataIn_1_payload_address_20;
    _zz_io_dataIn_1_payload_address_22 <= _zz_io_dataIn_1_payload_address_21;
    _zz_io_dataIn_1_payload_address_23 <= _zz_io_dataIn_1_payload_address_22;
    _zz_io_dataIn_1_payload_address_24 <= _zz_io_dataIn_1_payload_address_23;
    _zz_io_dataIn_1_payload_address_25 <= _zz_io_dataIn_1_payload_address_24;
    _zz_io_dataIn_1_payload_address_26 <= _zz_io_dataIn_1_payload_address_25;
    _zz_io_dataIn_1_payload_address_27 <= _zz_io_dataIn_1_payload_address_26;
    _zz_io_dataIn_1_payload_address_28 <= _zz_io_dataIn_1_payload_address_27;
    _zz_io_dataIn_1_payload_address_29 <= _zz_io_dataIn_1_payload_address_28;
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      _zz_io_dataIn_1_valid_35 <= 1'b0;
      _zz_io_dataIn_1_valid_36 <= 1'b0;
      _zz_io_dataIn_1_valid_37 <= 1'b0;
      _zz_io_dataIn_1_valid_38 <= 1'b0;
      _zz_io_dataIn_1_valid_39 <= 1'b0;
      _zz_io_dataIn_1_valid_40 <= 1'b0;
      _zz_io_dataIn_1_valid_41 <= 1'b0;
      _zz_io_dataIn_1_valid_42 <= 1'b0;
      _zz_io_dataIn_1_valid_43 <= 1'b0;
      _zz_io_dataIn_1_valid_44 <= 1'b0;
      _zz_io_dataIn_1_valid_45 <= 1'b0;
      _zz_io_dataIn_1_valid_46 <= 1'b0;
      _zz_io_dataIn_1_valid_47 <= 1'b0;
      _zz_io_dataIn_1_valid_48 <= 1'b0;
      _zz_io_dataIn_1_valid_49 <= 1'b0;
      _zz_io_dataIn_1_valid_50 <= 1'b0;
      _zz_io_dataIn_1_valid_51 <= 1'b0;
      _zz_io_dataIn_1_valid_52 <= 1'b0;
      _zz_io_dataIn_1_valid_53 <= 1'b0;
      _zz_io_dataIn_1_valid_54 <= 1'b0;
      _zz_io_dataIn_1_valid_55 <= 1'b0;
      _zz_io_dataIn_1_valid_56 <= 1'b0;
      _zz_io_dataIn_1_valid_57 <= 1'b0;
      _zz_io_dataIn_1_valid_58 <= 1'b0;
      _zz_io_dataIn_1_valid_59 <= 1'b0;
      _zz_io_dataIn_1_valid_60 <= 1'b0;
      _zz_io_dataIn_1_valid_61 <= 1'b0;
      _zz_io_dataIn_1_valid_62 <= 1'b0;
      _zz_io_dataIn_1_valid_63 <= 1'b0;
      _zz_io_dataIn_1_valid_64 <= 1'b0;
    end else begin
      _zz_io_dataIn_1_valid_35 <= (((fsm_stateReg & fsm_enumDef_stage2) != 4'b0000) && (! stage2_calCnt_value[1]));
      _zz_io_dataIn_1_valid_36 <= _zz_io_dataIn_1_valid_35;
      _zz_io_dataIn_1_valid_37 <= _zz_io_dataIn_1_valid_36;
      _zz_io_dataIn_1_valid_38 <= _zz_io_dataIn_1_valid_37;
      _zz_io_dataIn_1_valid_39 <= _zz_io_dataIn_1_valid_38;
      _zz_io_dataIn_1_valid_40 <= _zz_io_dataIn_1_valid_39;
      _zz_io_dataIn_1_valid_41 <= _zz_io_dataIn_1_valid_40;
      _zz_io_dataIn_1_valid_42 <= _zz_io_dataIn_1_valid_41;
      _zz_io_dataIn_1_valid_43 <= _zz_io_dataIn_1_valid_42;
      _zz_io_dataIn_1_valid_44 <= _zz_io_dataIn_1_valid_43;
      _zz_io_dataIn_1_valid_45 <= _zz_io_dataIn_1_valid_44;
      _zz_io_dataIn_1_valid_46 <= _zz_io_dataIn_1_valid_45;
      _zz_io_dataIn_1_valid_47 <= _zz_io_dataIn_1_valid_46;
      _zz_io_dataIn_1_valid_48 <= _zz_io_dataIn_1_valid_47;
      _zz_io_dataIn_1_valid_49 <= _zz_io_dataIn_1_valid_48;
      _zz_io_dataIn_1_valid_50 <= _zz_io_dataIn_1_valid_49;
      _zz_io_dataIn_1_valid_51 <= _zz_io_dataIn_1_valid_50;
      _zz_io_dataIn_1_valid_52 <= _zz_io_dataIn_1_valid_51;
      _zz_io_dataIn_1_valid_53 <= _zz_io_dataIn_1_valid_52;
      _zz_io_dataIn_1_valid_54 <= _zz_io_dataIn_1_valid_53;
      _zz_io_dataIn_1_valid_55 <= _zz_io_dataIn_1_valid_54;
      _zz_io_dataIn_1_valid_56 <= _zz_io_dataIn_1_valid_55;
      _zz_io_dataIn_1_valid_57 <= _zz_io_dataIn_1_valid_56;
      _zz_io_dataIn_1_valid_58 <= _zz_io_dataIn_1_valid_57;
      _zz_io_dataIn_1_valid_59 <= _zz_io_dataIn_1_valid_58;
      _zz_io_dataIn_1_valid_60 <= _zz_io_dataIn_1_valid_59;
      _zz_io_dataIn_1_valid_61 <= _zz_io_dataIn_1_valid_60;
      _zz_io_dataIn_1_valid_62 <= _zz_io_dataIn_1_valid_61;
      _zz_io_dataIn_1_valid_63 <= _zz_io_dataIn_1_valid_62;
      _zz_io_dataIn_1_valid_64 <= _zz_io_dataIn_1_valid_63;
    end
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      _zz_io_dataIn_1_valid_65 <= 1'b0;
      _zz_io_dataIn_1_valid_66 <= 1'b0;
      _zz_io_dataIn_1_valid_67 <= 1'b0;
      _zz_io_dataIn_1_valid_68 <= 1'b0;
      _zz_io_dataIn_1_valid_69 <= 1'b0;
      _zz_io_dataIn_1_valid_70 <= 1'b0;
      _zz_io_dataIn_1_valid_71 <= 1'b0;
      _zz_io_dataIn_1_valid_72 <= 1'b0;
      _zz_io_dataIn_1_valid_73 <= 1'b0;
      _zz_io_dataIn_1_valid_74 <= 1'b0;
      _zz_io_dataIn_1_valid_75 <= 1'b0;
      _zz_io_dataIn_1_valid_76 <= 1'b0;
      _zz_io_dataIn_1_valid_77 <= 1'b0;
      _zz_io_dataIn_1_valid_78 <= 1'b0;
      _zz_io_dataIn_1_valid_79 <= 1'b0;
      _zz_io_dataIn_1_valid_80 <= 1'b0;
      _zz_io_dataIn_1_valid_81 <= 1'b0;
      _zz_io_dataIn_1_valid_82 <= 1'b0;
      _zz_io_dataIn_1_valid_83 <= 1'b0;
      _zz_io_dataIn_1_valid_84 <= 1'b0;
      _zz_io_dataIn_1_valid_85 <= 1'b0;
      _zz_io_dataIn_1_valid_86 <= 1'b0;
      _zz_io_dataIn_1_valid_87 <= 1'b0;
      _zz_io_dataIn_1_valid_88 <= 1'b0;
      _zz_io_dataIn_1_valid_89 <= 1'b0;
      _zz_io_dataIn_1_valid_90 <= 1'b0;
      _zz_io_dataIn_1_valid_91 <= 1'b0;
      _zz_io_dataIn_1_valid_92 <= 1'b0;
      _zz_io_dataIn_1_valid_93 <= 1'b0;
      _zz_io_dataIn_1_valid_94 <= 1'b0;
    end else begin
      _zz_io_dataIn_1_valid_65 <= ((stage3_doubleWaitCnt_value == 9'h001) || (stage3_addWaitCnt_value == 9'h001));
      _zz_io_dataIn_1_valid_66 <= _zz_io_dataIn_1_valid_65;
      _zz_io_dataIn_1_valid_67 <= _zz_io_dataIn_1_valid_66;
      _zz_io_dataIn_1_valid_68 <= _zz_io_dataIn_1_valid_67;
      _zz_io_dataIn_1_valid_69 <= _zz_io_dataIn_1_valid_68;
      _zz_io_dataIn_1_valid_70 <= _zz_io_dataIn_1_valid_69;
      _zz_io_dataIn_1_valid_71 <= _zz_io_dataIn_1_valid_70;
      _zz_io_dataIn_1_valid_72 <= _zz_io_dataIn_1_valid_71;
      _zz_io_dataIn_1_valid_73 <= _zz_io_dataIn_1_valid_72;
      _zz_io_dataIn_1_valid_74 <= _zz_io_dataIn_1_valid_73;
      _zz_io_dataIn_1_valid_75 <= _zz_io_dataIn_1_valid_74;
      _zz_io_dataIn_1_valid_76 <= _zz_io_dataIn_1_valid_75;
      _zz_io_dataIn_1_valid_77 <= _zz_io_dataIn_1_valid_76;
      _zz_io_dataIn_1_valid_78 <= _zz_io_dataIn_1_valid_77;
      _zz_io_dataIn_1_valid_79 <= _zz_io_dataIn_1_valid_78;
      _zz_io_dataIn_1_valid_80 <= _zz_io_dataIn_1_valid_79;
      _zz_io_dataIn_1_valid_81 <= _zz_io_dataIn_1_valid_80;
      _zz_io_dataIn_1_valid_82 <= _zz_io_dataIn_1_valid_81;
      _zz_io_dataIn_1_valid_83 <= _zz_io_dataIn_1_valid_82;
      _zz_io_dataIn_1_valid_84 <= _zz_io_dataIn_1_valid_83;
      _zz_io_dataIn_1_valid_85 <= _zz_io_dataIn_1_valid_84;
      _zz_io_dataIn_1_valid_86 <= _zz_io_dataIn_1_valid_85;
      _zz_io_dataIn_1_valid_87 <= _zz_io_dataIn_1_valid_86;
      _zz_io_dataIn_1_valid_88 <= _zz_io_dataIn_1_valid_87;
      _zz_io_dataIn_1_valid_89 <= _zz_io_dataIn_1_valid_88;
      _zz_io_dataIn_1_valid_90 <= _zz_io_dataIn_1_valid_89;
      _zz_io_dataIn_1_valid_91 <= _zz_io_dataIn_1_valid_90;
      _zz_io_dataIn_1_valid_92 <= _zz_io_dataIn_1_valid_91;
      _zz_io_dataIn_1_valid_93 <= _zz_io_dataIn_1_valid_92;
      _zz_io_dataIn_1_valid_94 <= _zz_io_dataIn_1_valid_93;
    end
  end

  always @(posedge clk) begin
    pippenger_1_dataRam_0_io_rData_1_regNext_X_1 <= dataRam_0_io_rData_1_X;
    pippenger_1_dataRam_0_io_rData_1_regNext_Y_1 <= dataRam_0_io_rData_1_Y;
    pippenger_1_dataRam_0_io_rData_1_regNext_Z_1 <= dataRam_0_io_rData_1_Z;
    pippenger_1_dataRam_0_io_rData_1_regNext_T_1 <= dataRam_0_io_rData_1_T;
    _zz_io_dataIn_1_payload_address_30 <= (stage3_GCnt_value - _zz__zz_io_dataIn_1_payload_address_30);
    _zz_io_dataIn_1_payload_address_31 <= _zz_io_dataIn_1_payload_address_30;
    _zz_io_dataIn_1_payload_address_32 <= _zz_io_dataIn_1_payload_address_31;
    _zz_io_dataIn_1_payload_address_33 <= _zz_io_dataIn_1_payload_address_32;
    _zz_io_dataIn_1_payload_address_34 <= _zz_io_dataIn_1_payload_address_33;
    _zz_io_dataIn_1_payload_address_35 <= _zz_io_dataIn_1_payload_address_34;
    _zz_io_dataIn_1_payload_address_36 <= _zz_io_dataIn_1_payload_address_35;
    _zz_io_dataIn_1_payload_address_37 <= _zz_io_dataIn_1_payload_address_36;
    _zz_io_dataIn_1_payload_address_38 <= _zz_io_dataIn_1_payload_address_37;
    _zz_io_dataIn_1_payload_address_39 <= _zz_io_dataIn_1_payload_address_38;
    _zz_io_dataIn_1_payload_address_40 <= _zz_io_dataIn_1_payload_address_39;
    _zz_io_dataIn_1_payload_address_41 <= _zz_io_dataIn_1_payload_address_40;
    _zz_io_dataIn_1_payload_address_42 <= _zz_io_dataIn_1_payload_address_41;
    _zz_io_dataIn_1_payload_address_43 <= _zz_io_dataIn_1_payload_address_42;
    _zz_io_dataIn_1_payload_address_44 <= _zz_io_dataIn_1_payload_address_43;
    _zz_io_dataIn_1_payload_address_45 <= _zz_io_dataIn_1_payload_address_44;
    _zz_io_dataIn_1_payload_address_46 <= _zz_io_dataIn_1_payload_address_45;
    _zz_io_dataIn_1_payload_address_47 <= _zz_io_dataIn_1_payload_address_46;
    _zz_io_dataIn_1_payload_address_48 <= _zz_io_dataIn_1_payload_address_47;
    _zz_io_dataIn_1_payload_address_49 <= _zz_io_dataIn_1_payload_address_48;
    _zz_io_dataIn_1_payload_address_50 <= _zz_io_dataIn_1_payload_address_49;
    _zz_io_dataIn_1_payload_address_51 <= _zz_io_dataIn_1_payload_address_50;
    _zz_io_dataIn_1_payload_address_52 <= _zz_io_dataIn_1_payload_address_51;
    _zz_io_dataIn_1_payload_address_53 <= _zz_io_dataIn_1_payload_address_52;
    _zz_io_dataIn_1_payload_address_54 <= _zz_io_dataIn_1_payload_address_53;
    _zz_io_dataIn_1_payload_address_55 <= _zz_io_dataIn_1_payload_address_54;
    _zz_io_dataIn_1_payload_address_56 <= _zz_io_dataIn_1_payload_address_55;
    _zz_io_dataIn_1_payload_address_57 <= _zz_io_dataIn_1_payload_address_56;
    _zz_io_dataIn_1_payload_address_58 <= _zz_io_dataIn_1_payload_address_57;
    _zz_io_dataIn_1_payload_address_59 <= _zz_io_dataIn_1_payload_address_58;
  end


endmodule

module PNeg (
  input      [376:0]  io_a_X,
  input      [376:0]  io_a_Y,
  input      [376:0]  io_a_Z,
  input      [376:0]  io_a_T,
  output     [376:0]  io_n_X,
  output     [376:0]  io_n_Y,
  output     [376:0]  io_n_Z,
  output     [376:0]  io_n_T,
  input               clk,
  input               resetn
);

  wire       [377:0]  sub_io_s;
  reg        [376:0]  io_a_X_delay_1;
  reg        [376:0]  io_a_X_delay_2;
  reg        [376:0]  io_a_X_delay_3;
  reg        [376:0]  io_a_X_delay_4;
  reg        [376:0]  io_a_X_delay_5;
  reg        [376:0]  io_a_X_delay_6;
  reg        [376:0]  io_a_T_delay_1;
  reg        [376:0]  io_a_T_delay_2;
  reg        [376:0]  io_a_T_delay_3;
  reg        [376:0]  io_a_T_delay_4;
  reg        [376:0]  io_a_T_delay_5;
  reg        [376:0]  io_a_T_delay_6;

  BADD sub (
    .io_a   (377'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001), //i
    .io_b   (io_a_Y[376:0]                                                                                       ), //i
    .io_c   (1'b1                                                                                                ), //i
    .io_s   (sub_io_s[377:0]                                                                                     ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  assign io_n_X = io_a_X_delay_6;
  assign io_n_Y = sub_io_s[376:0];
  assign io_n_Z = 377'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000000;
  assign io_n_T = io_a_T_delay_6;
  always @(posedge clk) begin
    io_a_X_delay_1 <= io_a_X;
    io_a_X_delay_2 <= io_a_X_delay_1;
    io_a_X_delay_3 <= io_a_X_delay_2;
    io_a_X_delay_4 <= io_a_X_delay_3;
    io_a_X_delay_5 <= io_a_X_delay_4;
    io_a_X_delay_6 <= io_a_X_delay_5;
    io_a_T_delay_1 <= io_a_T;
    io_a_T_delay_2 <= io_a_T_delay_1;
    io_a_T_delay_3 <= io_a_T_delay_2;
    io_a_T_delay_4 <= io_a_T_delay_3;
    io_a_T_delay_5 <= io_a_T_delay_4;
    io_a_T_delay_6 <= io_a_T_delay_5;
  end


endmodule

module PAdd (
  input      [376:0]  io_a_X,
  input      [376:0]  io_a_Y,
  input      [376:0]  io_a_Z,
  input      [376:0]  io_a_T,
  input      [376:0]  io_b_X,
  input      [376:0]  io_b_Y,
  input      [376:0]  io_b_Z,
  input      [376:0]  io_b_T,
  output     [376:0]  io_s_X,
  output     [376:0]  io_s_Y,
  output     [376:0]  io_s_Z,
  output     [376:0]  io_s_T,
  input               clk,
  input               resetn
);

  wire       [377:0]  reduction_io_a;
  wire       [376:0]  mul_0_io_p;
  wire       [376:0]  mul_1_io_p;
  wire       [376:0]  mul_2_io_p;
  wire       [376:0]  mul_3_io_p;
  wire       [376:0]  mul_4_io_p;
  wire       [376:0]  mul_5_io_p;
  wire       [376:0]  mul_6_io_p;
  wire       [376:0]  mul_7_io_p;
  wire       [376:0]  cMul_io_p;
  wire       [376:0]  add_0_io_s;
  wire       [376:0]  add_1_io_s;
  wire       [376:0]  add_2_io_s;
  wire       [376:0]  add_3_io_s;
  wire       [376:0]  sub_0_io_s;
  wire       [376:0]  sub_1_io_s;
  wire       [376:0]  sub_2_io_s;
  wire       [376:0]  sub_3_io_s;
  wire       [376:0]  reduction_io_r;
  reg        [376:0]  io_a_T_delay_1;
  reg        [376:0]  io_a_T_delay_2;
  reg        [376:0]  io_a_T_delay_3;
  reg        [376:0]  io_a_T_delay_4;
  reg        [376:0]  io_a_T_delay_5;
  reg        [376:0]  io_a_T_delay_6;
  reg        [376:0]  io_a_T_delay_7;
  reg        [376:0]  io_a_T_delay_8;
  reg        [376:0]  io_a_T_delay_9;
  reg        [376:0]  io_a_T_delay_10;
  reg        [376:0]  io_a_T_delay_11;
  reg        [376:0]  io_a_T_delay_12;
  reg        [376:0]  io_a_T_delay_13;
  reg        [376:0]  io_a_T_delay_14;
  reg        [376:0]  io_a_T_delay_15;
  reg        [376:0]  io_a_T_delay_16;
  reg        [376:0]  io_a_T_delay_17;
  reg        [376:0]  io_a_T_delay_18;
  reg        [376:0]  io_a_T_delay_19;
  reg        [376:0]  io_a_T_delay_20;
  reg        [376:0]  io_a_T_delay_21;
  reg        [376:0]  io_a_T_delay_22;
  reg        [376:0]  io_a_T_delay_23;
  reg        [376:0]  io_a_T_delay_24;
  reg        [376:0]  io_a_T_delay_25;
  reg        [376:0]  io_a_T_delay_26;
  reg        [376:0]  io_a_T_delay_27;
  reg        [376:0]  io_a_T_delay_28;
  reg        [376:0]  io_a_T_delay_29;
  reg        [376:0]  io_a_T_delay_30;
  reg        [376:0]  io_a_T_delay_31;
  reg        [376:0]  io_a_T_delay_32;
  reg        [376:0]  io_a_T_delay_33;
  reg        [376:0]  io_a_T_delay_34;
  reg        [376:0]  io_a_T_delay_35;
  reg        [376:0]  io_a_T_delay_36;
  reg        [376:0]  io_a_T_delay_37;
  reg        [376:0]  io_a_T_delay_38;
  reg        [376:0]  io_a_T_delay_39;
  reg        [376:0]  io_a_T_delay_40;
  reg        [376:0]  io_a_T_delay_41;
  reg        [376:0]  io_a_T_delay_42;
  reg        [376:0]  io_a_T_delay_43;
  reg        [376:0]  io_a_T_delay_44;
  reg        [376:0]  io_a_T_delay_45;
  reg        [376:0]  io_a_T_delay_46;
  reg        [376:0]  io_a_T_delay_47;
  reg        [376:0]  io_a_T_delay_48;
  reg        [376:0]  io_a_T_delay_49;
  reg        [376:0]  io_a_T_delay_50;
  reg        [376:0]  io_a_T_delay_51;
  reg        [376:0]  io_a_T_delay_52;
  reg        [376:0]  io_a_T_delay_53;
  reg        [376:0]  io_a_T_delay_54;
  reg        [376:0]  io_a_T_delay_55;
  reg        [376:0]  io_a_T_delay_56;
  reg        [376:0]  io_a_T_delay_57;
  reg        [376:0]  io_a_T_delay_58;
  reg        [376:0]  io_a_T_delay_59;
  reg        [376:0]  io_a_T_delay_60;
  reg        [376:0]  io_a_T_delay_61;
  reg        [376:0]  io_a_T_delay_62;
  reg        [376:0]  io_a_T_delay_63;
  reg        [376:0]  io_a_T_delay_64;
  reg        [376:0]  io_a_T_delay_65;
  reg        [376:0]  io_a_T_delay_66;
  reg        [376:0]  io_a_T_delay_67;
  reg        [376:0]  io_a_T_delay_68;
  reg        [376:0]  io_a_T_delay_69;
  reg        [376:0]  io_a_T_delay_70;
  reg        [376:0]  io_a_T_delay_71;
  reg        [376:0]  io_a_T_delay_72;
  reg        [376:0]  io_a_T_delay_73;
  reg        [376:0]  io_a_T_delay_74;
  reg        [376:0]  io_a_T_delay_75;
  reg        [376:0]  io_a_T_delay_76;
  reg        [376:0]  io_a_T_delay_77;
  reg        [376:0]  io_a_T_delay_78;
  reg        [376:0]  io_a_T_delay_79;
  reg        [376:0]  io_a_T_delay_80;
  reg        [376:0]  io_a_T_delay_81;
  reg        [376:0]  io_a_T_delay_82;
  reg        [376:0]  io_a_T_delay_83;
  reg        [376:0]  io_a_T_delay_84;
  reg        [376:0]  adder_0_reduction_io_r_delay_1;
  reg        [376:0]  adder_0_reduction_io_r_delay_2;
  reg        [376:0]  adder_0_reduction_io_r_delay_3;
  reg        [376:0]  adder_0_reduction_io_r_delay_4;
  reg        [376:0]  adder_0_reduction_io_r_delay_5;
  reg        [376:0]  adder_0_reduction_io_r_delay_6;
  reg        [376:0]  adder_0_reduction_io_r_delay_7;
  reg        [376:0]  adder_0_reduction_io_r_delay_8;
  reg        [376:0]  adder_0_reduction_io_r_delay_9;
  reg        [376:0]  adder_0_reduction_io_r_delay_10;
  reg        [376:0]  adder_0_reduction_io_r_delay_11;
  reg        [376:0]  adder_0_reduction_io_r_delay_12;
  reg        [376:0]  adder_0_reduction_io_r_delay_13;
  reg        [376:0]  adder_0_reduction_io_r_delay_14;
  reg        [376:0]  adder_0_reduction_io_r_delay_15;
  reg        [376:0]  adder_0_reduction_io_r_delay_16;
  reg        [376:0]  adder_0_reduction_io_r_delay_17;
  reg        [376:0]  adder_0_reduction_io_r_delay_18;
  reg        [376:0]  adder_0_reduction_io_r_delay_19;
  reg        [376:0]  adder_0_reduction_io_r_delay_20;
  reg        [376:0]  adder_0_reduction_io_r_delay_21;
  reg        [376:0]  adder_0_reduction_io_r_delay_22;
  reg        [376:0]  adder_0_reduction_io_r_delay_23;
  reg        [376:0]  adder_0_reduction_io_r_delay_24;
  reg        [376:0]  adder_0_reduction_io_r_delay_25;
  reg        [376:0]  adder_0_reduction_io_r_delay_26;
  reg        [376:0]  adder_0_reduction_io_r_delay_27;
  reg        [376:0]  adder_0_reduction_io_r_delay_28;
  reg        [376:0]  adder_0_reduction_io_r_delay_29;
  reg        [376:0]  adder_0_reduction_io_r_delay_30;
  reg        [376:0]  adder_0_reduction_io_r_delay_31;
  reg        [376:0]  adder_0_reduction_io_r_delay_32;
  reg        [376:0]  adder_0_reduction_io_r_delay_33;
  reg        [376:0]  adder_0_reduction_io_r_delay_34;
  reg        [376:0]  adder_0_reduction_io_r_delay_35;
  reg        [376:0]  adder_0_reduction_io_r_delay_36;
  reg        [376:0]  adder_0_reduction_io_r_delay_37;
  reg        [376:0]  adder_0_reduction_io_r_delay_38;
  reg        [376:0]  adder_0_reduction_io_r_delay_39;
  reg        [376:0]  adder_0_reduction_io_r_delay_40;
  reg        [376:0]  adder_0_reduction_io_r_delay_41;
  reg        [376:0]  adder_0_reduction_io_r_delay_42;
  reg        [376:0]  adder_0_reduction_io_r_delay_43;
  reg        [376:0]  adder_0_reduction_io_r_delay_44;
  reg        [376:0]  adder_0_reduction_io_r_delay_45;
  reg        [376:0]  adder_0_reduction_io_r_delay_46;
  reg        [376:0]  adder_0_reduction_io_r_delay_47;
  reg        [376:0]  adder_0_reduction_io_r_delay_48;
  reg        [376:0]  adder_0_reduction_io_r_delay_49;
  reg        [376:0]  adder_0_reduction_io_r_delay_50;
  reg        [376:0]  adder_0_reduction_io_r_delay_51;
  reg        [376:0]  adder_0_reduction_io_r_delay_52;
  reg        [376:0]  adder_0_reduction_io_r_delay_53;
  reg        [376:0]  adder_0_reduction_io_r_delay_54;
  reg        [376:0]  adder_0_reduction_io_r_delay_55;
  reg        [376:0]  adder_0_reduction_io_r_delay_56;
  reg        [376:0]  adder_0_reduction_io_r_delay_57;
  reg        [376:0]  adder_0_reduction_io_r_delay_58;
  reg        [376:0]  adder_0_reduction_io_r_delay_59;
  reg        [376:0]  adder_0_reduction_io_r_delay_60;
  reg        [376:0]  adder_0_reduction_io_r_delay_61;
  reg        [376:0]  adder_0_reduction_io_r_delay_62;
  reg        [376:0]  adder_0_reduction_io_r_delay_63;
  reg        [376:0]  adder_0_reduction_io_r_delay_64;
  reg        [376:0]  adder_0_reduction_io_r_delay_65;
  reg        [376:0]  adder_0_reduction_io_r_delay_66;
  reg        [376:0]  adder_0_reduction_io_r_delay_67;
  reg        [376:0]  adder_0_reduction_io_r_delay_68;
  reg        [376:0]  adder_0_reduction_io_r_delay_69;
  reg        [376:0]  adder_0_reduction_io_r_delay_70;
  reg        [376:0]  adder_0_reduction_io_r_delay_71;
  reg        [376:0]  adder_0_reduction_io_r_delay_72;
  reg        [376:0]  adder_0_reduction_io_r_delay_73;
  reg        [376:0]  adder_0_reduction_io_r_delay_74;
  reg        [376:0]  adder_0_reduction_io_r_delay_75;
  reg        [376:0]  adder_0_reduction_io_r_delay_76;
  reg        [376:0]  R8;
  reg        [376:0]  adder_0_sub_2_io_s_delay_1;
  reg        [376:0]  adder_0_sub_2_io_s_delay_2;
  reg        [376:0]  adder_0_sub_2_io_s_delay_3;
  reg        [376:0]  adder_0_sub_2_io_s_delay_4;
  reg        [376:0]  adder_0_sub_2_io_s_delay_5;
  reg        [376:0]  adder_0_sub_2_io_s_delay_6;
  reg        [376:0]  adder_0_sub_2_io_s_delay_7;
  reg        [376:0]  adder_0_sub_2_io_s_delay_8;
  reg        [376:0]  adder_0_sub_2_io_s_delay_9;
  reg        [376:0]  adder_0_sub_2_io_s_delay_10;
  reg        [376:0]  adder_0_sub_2_io_s_delay_11;
  reg        [376:0]  adder_0_sub_2_io_s_delay_12;
  reg        [376:0]  adder_0_sub_2_io_s_delay_13;
  reg        [376:0]  adder_0_sub_2_io_s_delay_14;
  reg        [376:0]  adder_0_sub_2_io_s_delay_15;
  reg        [376:0]  adder_0_sub_2_io_s_delay_16;
  reg        [376:0]  adder_0_sub_2_io_s_delay_17;
  reg        [376:0]  adder_0_sub_2_io_s_delay_18;
  reg        [376:0]  adder_0_sub_2_io_s_delay_19;
  reg        [376:0]  adder_0_sub_2_io_s_delay_20;
  reg        [376:0]  adder_0_sub_2_io_s_delay_21;
  reg        [376:0]  adder_0_sub_2_io_s_delay_22;
  reg        [376:0]  adder_0_sub_2_io_s_delay_23;
  reg        [376:0]  adder_0_sub_2_io_s_delay_24;
  reg        [376:0]  adder_0_sub_2_io_s_delay_25;
  reg        [376:0]  adder_0_sub_2_io_s_delay_26;
  reg        [376:0]  adder_0_sub_2_io_s_delay_27;
  reg        [376:0]  adder_0_sub_2_io_s_delay_28;
  reg        [376:0]  adder_0_sub_2_io_s_delay_29;
  reg        [376:0]  adder_0_sub_2_io_s_delay_30;
  reg        [376:0]  adder_0_sub_2_io_s_delay_31;
  reg        [376:0]  adder_0_sub_2_io_s_delay_32;
  reg        [376:0]  adder_0_sub_2_io_s_delay_33;
  reg        [376:0]  adder_0_sub_2_io_s_delay_34;
  reg        [376:0]  adder_0_sub_2_io_s_delay_35;
  reg        [376:0]  adder_0_sub_2_io_s_delay_36;
  reg        [376:0]  adder_0_sub_2_io_s_delay_37;
  reg        [376:0]  adder_0_sub_2_io_s_delay_38;
  reg        [376:0]  adder_0_sub_2_io_s_delay_39;
  reg        [376:0]  adder_0_sub_2_io_s_delay_40;
  reg        [376:0]  adder_0_sub_2_io_s_delay_41;
  reg        [376:0]  adder_0_sub_2_io_s_delay_42;
  reg        [376:0]  adder_0_sub_2_io_s_delay_43;
  reg        [376:0]  adder_0_sub_2_io_s_delay_44;
  reg        [376:0]  adder_0_sub_2_io_s_delay_45;
  reg        [376:0]  adder_0_sub_2_io_s_delay_46;
  reg        [376:0]  adder_0_sub_2_io_s_delay_47;
  reg        [376:0]  adder_0_sub_2_io_s_delay_48;
  reg        [376:0]  adder_0_sub_2_io_s_delay_49;
  reg        [376:0]  adder_0_sub_2_io_s_delay_50;
  reg        [376:0]  adder_0_sub_2_io_s_delay_51;
  reg        [376:0]  adder_0_sub_2_io_s_delay_52;
  reg        [376:0]  adder_0_sub_2_io_s_delay_53;
  reg        [376:0]  adder_0_sub_2_io_s_delay_54;
  reg        [376:0]  adder_0_sub_2_io_s_delay_55;
  reg        [376:0]  adder_0_sub_2_io_s_delay_56;
  reg        [376:0]  adder_0_sub_2_io_s_delay_57;
  reg        [376:0]  adder_0_sub_2_io_s_delay_58;
  reg        [376:0]  adder_0_sub_2_io_s_delay_59;
  reg        [376:0]  adder_0_sub_2_io_s_delay_60;
  reg        [376:0]  adder_0_sub_2_io_s_delay_61;
  reg        [376:0]  adder_0_sub_2_io_s_delay_62;
  reg        [376:0]  adder_0_sub_2_io_s_delay_63;
  reg        [376:0]  adder_0_sub_2_io_s_delay_64;
  reg        [376:0]  adder_0_sub_2_io_s_delay_65;
  reg        [376:0]  adder_0_sub_2_io_s_delay_66;
  reg        [376:0]  adder_0_sub_2_io_s_delay_67;
  reg        [376:0]  adder_0_sub_2_io_s_delay_68;
  reg        [376:0]  adder_0_sub_2_io_s_delay_69;
  reg        [376:0]  adder_0_sub_2_io_s_delay_70;
  reg        [376:0]  adder_0_sub_2_io_s_delay_71;
  reg        [376:0]  adder_0_sub_2_io_s_delay_72;
  reg        [376:0]  adder_0_sub_2_io_s_delay_73;
  reg        [376:0]  adder_0_sub_2_io_s_delay_74;
  reg        [376:0]  adder_0_sub_2_io_s_delay_75;
  reg        [376:0]  R9;
  reg        [376:0]  adder_0_add_3_io_s_delay_1;
  reg        [376:0]  adder_0_add_3_io_s_delay_2;
  reg        [376:0]  adder_0_add_3_io_s_delay_3;
  reg        [376:0]  adder_0_add_3_io_s_delay_4;
  reg        [376:0]  adder_0_add_3_io_s_delay_5;
  reg        [376:0]  adder_0_add_3_io_s_delay_6;
  reg        [376:0]  adder_0_add_3_io_s_delay_7;
  reg        [376:0]  adder_0_add_3_io_s_delay_8;
  reg        [376:0]  adder_0_add_3_io_s_delay_9;
  reg        [376:0]  adder_0_add_3_io_s_delay_10;
  reg        [376:0]  adder_0_add_3_io_s_delay_11;
  reg        [376:0]  adder_0_add_3_io_s_delay_12;
  reg        [376:0]  adder_0_add_3_io_s_delay_13;
  reg        [376:0]  adder_0_add_3_io_s_delay_14;
  reg        [376:0]  adder_0_add_3_io_s_delay_15;
  reg        [376:0]  adder_0_add_3_io_s_delay_16;
  reg        [376:0]  adder_0_add_3_io_s_delay_17;
  reg        [376:0]  adder_0_add_3_io_s_delay_18;
  reg        [376:0]  adder_0_add_3_io_s_delay_19;
  reg        [376:0]  adder_0_add_3_io_s_delay_20;
  reg        [376:0]  adder_0_add_3_io_s_delay_21;
  reg        [376:0]  adder_0_add_3_io_s_delay_22;
  reg        [376:0]  adder_0_add_3_io_s_delay_23;
  reg        [376:0]  adder_0_add_3_io_s_delay_24;
  reg        [376:0]  adder_0_add_3_io_s_delay_25;
  reg        [376:0]  adder_0_add_3_io_s_delay_26;
  reg        [376:0]  adder_0_add_3_io_s_delay_27;
  reg        [376:0]  adder_0_add_3_io_s_delay_28;
  reg        [376:0]  adder_0_add_3_io_s_delay_29;
  reg        [376:0]  adder_0_add_3_io_s_delay_30;
  reg        [376:0]  adder_0_add_3_io_s_delay_31;
  reg        [376:0]  adder_0_add_3_io_s_delay_32;
  reg        [376:0]  adder_0_add_3_io_s_delay_33;
  reg        [376:0]  adder_0_add_3_io_s_delay_34;
  reg        [376:0]  adder_0_add_3_io_s_delay_35;
  reg        [376:0]  adder_0_add_3_io_s_delay_36;
  reg        [376:0]  adder_0_add_3_io_s_delay_37;
  reg        [376:0]  adder_0_add_3_io_s_delay_38;
  reg        [376:0]  adder_0_add_3_io_s_delay_39;
  reg        [376:0]  adder_0_add_3_io_s_delay_40;
  reg        [376:0]  adder_0_add_3_io_s_delay_41;
  reg        [376:0]  adder_0_add_3_io_s_delay_42;
  reg        [376:0]  adder_0_add_3_io_s_delay_43;
  reg        [376:0]  adder_0_add_3_io_s_delay_44;
  reg        [376:0]  adder_0_add_3_io_s_delay_45;
  reg        [376:0]  adder_0_add_3_io_s_delay_46;
  reg        [376:0]  adder_0_add_3_io_s_delay_47;
  reg        [376:0]  adder_0_add_3_io_s_delay_48;
  reg        [376:0]  adder_0_add_3_io_s_delay_49;
  reg        [376:0]  adder_0_add_3_io_s_delay_50;
  reg        [376:0]  adder_0_add_3_io_s_delay_51;
  reg        [376:0]  adder_0_add_3_io_s_delay_52;
  reg        [376:0]  adder_0_add_3_io_s_delay_53;
  reg        [376:0]  adder_0_add_3_io_s_delay_54;
  reg        [376:0]  adder_0_add_3_io_s_delay_55;
  reg        [376:0]  adder_0_add_3_io_s_delay_56;
  reg        [376:0]  adder_0_add_3_io_s_delay_57;
  reg        [376:0]  adder_0_add_3_io_s_delay_58;
  reg        [376:0]  adder_0_add_3_io_s_delay_59;
  reg        [376:0]  adder_0_add_3_io_s_delay_60;
  reg        [376:0]  adder_0_add_3_io_s_delay_61;
  reg        [376:0]  adder_0_add_3_io_s_delay_62;
  reg        [376:0]  adder_0_add_3_io_s_delay_63;
  reg        [376:0]  adder_0_add_3_io_s_delay_64;
  reg        [376:0]  adder_0_add_3_io_s_delay_65;
  reg        [376:0]  adder_0_add_3_io_s_delay_66;
  reg        [376:0]  adder_0_add_3_io_s_delay_67;
  reg        [376:0]  adder_0_add_3_io_s_delay_68;
  reg        [376:0]  adder_0_add_3_io_s_delay_69;
  reg        [376:0]  adder_0_add_3_io_s_delay_70;
  reg        [376:0]  adder_0_add_3_io_s_delay_71;
  reg        [376:0]  adder_0_add_3_io_s_delay_72;
  reg        [376:0]  adder_0_add_3_io_s_delay_73;
  reg        [376:0]  adder_0_add_3_io_s_delay_74;
  reg        [376:0]  adder_0_add_3_io_s_delay_75;
  reg        [376:0]  R12;

  KaratsubaMMUL mul_0 (
    .io_a   (sub_0_io_s[376:0]), //i
    .io_b   (sub_1_io_s[376:0]), //i
    .io_p   (mul_0_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL mul_1 (
    .io_a   (add_0_io_s[376:0]), //i
    .io_b   (add_1_io_s[376:0]), //i
    .io_p   (mul_1_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL mul_2 (
    .io_a   (io_a_T_delay_84[376:0]), //i
    .io_b   (cMul_io_p[376:0]      ), //i
    .io_p   (mul_2_io_p[376:0]     ), //o
    .clk    (clk                   ), //i
    .resetn (resetn                )  //i
  );
  KaratsubaMMUL mul_3 (
    .io_a   (io_a_Z[376:0]    ), //i
    .io_b   (io_b_Z[376:0]    ), //i
    .io_p   (mul_3_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL mul_4 (
    .io_a   (R9[376:0]        ), //i
    .io_b   (sub_3_io_s[376:0]), //i
    .io_p   (mul_4_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL mul_5 (
    .io_a   (add_2_io_s[376:0]), //i
    .io_b   (R12[376:0]       ), //i
    .io_p   (mul_5_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL mul_6 (
    .io_a   (sub_3_io_s[376:0]), //i
    .io_b   (add_2_io_s[376:0]), //i
    .io_p   (mul_6_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL mul_7 (
    .io_a   (R9[376:0]        ), //i
    .io_b   (R12[376:0]       ), //i
    .io_p   (mul_7_io_p[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  KaratsubaMMUL cMul (
    .io_a   (io_b_T[376:0]                                                                                       ), //i
    .io_b   (377'h196bab03169a4f2ca0b7670ae65fc7437786998c1a32d217f165b2fe0b32139735d947870e3d3e4e02c125684d6e016), //i
    .io_p   (cMul_io_p[376:0]                                                                                    ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  MADD add_0 (
    .io_a   (io_a_Y[376:0]    ), //i
    .io_b   (io_a_X[376:0]    ), //i
    .io_s   (add_0_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD add_1 (
    .io_a   (io_b_Y[376:0]    ), //i
    .io_b   (io_b_X[376:0]    ), //i
    .io_s   (add_1_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD add_2 (
    .io_a   (R8[376:0]        ), //i
    .io_b   (mul_2_io_p[376:0]), //i
    .io_s   (add_2_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD add_3 (
    .io_a   (mul_1_io_p[376:0]), //i
    .io_b   (mul_0_io_p[376:0]), //i
    .io_s   (add_3_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_4 sub_0 (
    .io_a   (io_a_Y[376:0]    ), //i
    .io_b   (io_a_X[376:0]    ), //i
    .io_s   (sub_0_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_4 sub_1 (
    .io_a   (io_b_Y[376:0]    ), //i
    .io_b   (io_b_X[376:0]    ), //i
    .io_s   (sub_1_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_4 sub_2 (
    .io_a   (mul_1_io_p[376:0]), //i
    .io_b   (mul_0_io_p[376:0]), //i
    .io_s   (sub_2_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  MADD_4 sub_3 (
    .io_a   (R8[376:0]        ), //i
    .io_b   (mul_2_io_p[376:0]), //i
    .io_s   (sub_3_io_s[376:0]), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  FineReduction reduction (
    .io_a   (reduction_io_a[377:0]), //i
    .io_r   (reduction_io_r[376:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign reduction_io_a = ({1'd0,mul_3_io_p} <<< 1);
  assign io_s_X = mul_4_io_p;
  assign io_s_Y = mul_5_io_p;
  assign io_s_Z = mul_6_io_p;
  assign io_s_T = mul_7_io_p;
  always @(posedge clk) begin
    io_a_T_delay_1 <= io_a_T;
    io_a_T_delay_2 <= io_a_T_delay_1;
    io_a_T_delay_3 <= io_a_T_delay_2;
    io_a_T_delay_4 <= io_a_T_delay_3;
    io_a_T_delay_5 <= io_a_T_delay_4;
    io_a_T_delay_6 <= io_a_T_delay_5;
    io_a_T_delay_7 <= io_a_T_delay_6;
    io_a_T_delay_8 <= io_a_T_delay_7;
    io_a_T_delay_9 <= io_a_T_delay_8;
    io_a_T_delay_10 <= io_a_T_delay_9;
    io_a_T_delay_11 <= io_a_T_delay_10;
    io_a_T_delay_12 <= io_a_T_delay_11;
    io_a_T_delay_13 <= io_a_T_delay_12;
    io_a_T_delay_14 <= io_a_T_delay_13;
    io_a_T_delay_15 <= io_a_T_delay_14;
    io_a_T_delay_16 <= io_a_T_delay_15;
    io_a_T_delay_17 <= io_a_T_delay_16;
    io_a_T_delay_18 <= io_a_T_delay_17;
    io_a_T_delay_19 <= io_a_T_delay_18;
    io_a_T_delay_20 <= io_a_T_delay_19;
    io_a_T_delay_21 <= io_a_T_delay_20;
    io_a_T_delay_22 <= io_a_T_delay_21;
    io_a_T_delay_23 <= io_a_T_delay_22;
    io_a_T_delay_24 <= io_a_T_delay_23;
    io_a_T_delay_25 <= io_a_T_delay_24;
    io_a_T_delay_26 <= io_a_T_delay_25;
    io_a_T_delay_27 <= io_a_T_delay_26;
    io_a_T_delay_28 <= io_a_T_delay_27;
    io_a_T_delay_29 <= io_a_T_delay_28;
    io_a_T_delay_30 <= io_a_T_delay_29;
    io_a_T_delay_31 <= io_a_T_delay_30;
    io_a_T_delay_32 <= io_a_T_delay_31;
    io_a_T_delay_33 <= io_a_T_delay_32;
    io_a_T_delay_34 <= io_a_T_delay_33;
    io_a_T_delay_35 <= io_a_T_delay_34;
    io_a_T_delay_36 <= io_a_T_delay_35;
    io_a_T_delay_37 <= io_a_T_delay_36;
    io_a_T_delay_38 <= io_a_T_delay_37;
    io_a_T_delay_39 <= io_a_T_delay_38;
    io_a_T_delay_40 <= io_a_T_delay_39;
    io_a_T_delay_41 <= io_a_T_delay_40;
    io_a_T_delay_42 <= io_a_T_delay_41;
    io_a_T_delay_43 <= io_a_T_delay_42;
    io_a_T_delay_44 <= io_a_T_delay_43;
    io_a_T_delay_45 <= io_a_T_delay_44;
    io_a_T_delay_46 <= io_a_T_delay_45;
    io_a_T_delay_47 <= io_a_T_delay_46;
    io_a_T_delay_48 <= io_a_T_delay_47;
    io_a_T_delay_49 <= io_a_T_delay_48;
    io_a_T_delay_50 <= io_a_T_delay_49;
    io_a_T_delay_51 <= io_a_T_delay_50;
    io_a_T_delay_52 <= io_a_T_delay_51;
    io_a_T_delay_53 <= io_a_T_delay_52;
    io_a_T_delay_54 <= io_a_T_delay_53;
    io_a_T_delay_55 <= io_a_T_delay_54;
    io_a_T_delay_56 <= io_a_T_delay_55;
    io_a_T_delay_57 <= io_a_T_delay_56;
    io_a_T_delay_58 <= io_a_T_delay_57;
    io_a_T_delay_59 <= io_a_T_delay_58;
    io_a_T_delay_60 <= io_a_T_delay_59;
    io_a_T_delay_61 <= io_a_T_delay_60;
    io_a_T_delay_62 <= io_a_T_delay_61;
    io_a_T_delay_63 <= io_a_T_delay_62;
    io_a_T_delay_64 <= io_a_T_delay_63;
    io_a_T_delay_65 <= io_a_T_delay_64;
    io_a_T_delay_66 <= io_a_T_delay_65;
    io_a_T_delay_67 <= io_a_T_delay_66;
    io_a_T_delay_68 <= io_a_T_delay_67;
    io_a_T_delay_69 <= io_a_T_delay_68;
    io_a_T_delay_70 <= io_a_T_delay_69;
    io_a_T_delay_71 <= io_a_T_delay_70;
    io_a_T_delay_72 <= io_a_T_delay_71;
    io_a_T_delay_73 <= io_a_T_delay_72;
    io_a_T_delay_74 <= io_a_T_delay_73;
    io_a_T_delay_75 <= io_a_T_delay_74;
    io_a_T_delay_76 <= io_a_T_delay_75;
    io_a_T_delay_77 <= io_a_T_delay_76;
    io_a_T_delay_78 <= io_a_T_delay_77;
    io_a_T_delay_79 <= io_a_T_delay_78;
    io_a_T_delay_80 <= io_a_T_delay_79;
    io_a_T_delay_81 <= io_a_T_delay_80;
    io_a_T_delay_82 <= io_a_T_delay_81;
    io_a_T_delay_83 <= io_a_T_delay_82;
    io_a_T_delay_84 <= io_a_T_delay_83;
    adder_0_reduction_io_r_delay_1 <= reduction_io_r;
    adder_0_reduction_io_r_delay_2 <= adder_0_reduction_io_r_delay_1;
    adder_0_reduction_io_r_delay_3 <= adder_0_reduction_io_r_delay_2;
    adder_0_reduction_io_r_delay_4 <= adder_0_reduction_io_r_delay_3;
    adder_0_reduction_io_r_delay_5 <= adder_0_reduction_io_r_delay_4;
    adder_0_reduction_io_r_delay_6 <= adder_0_reduction_io_r_delay_5;
    adder_0_reduction_io_r_delay_7 <= adder_0_reduction_io_r_delay_6;
    adder_0_reduction_io_r_delay_8 <= adder_0_reduction_io_r_delay_7;
    adder_0_reduction_io_r_delay_9 <= adder_0_reduction_io_r_delay_8;
    adder_0_reduction_io_r_delay_10 <= adder_0_reduction_io_r_delay_9;
    adder_0_reduction_io_r_delay_11 <= adder_0_reduction_io_r_delay_10;
    adder_0_reduction_io_r_delay_12 <= adder_0_reduction_io_r_delay_11;
    adder_0_reduction_io_r_delay_13 <= adder_0_reduction_io_r_delay_12;
    adder_0_reduction_io_r_delay_14 <= adder_0_reduction_io_r_delay_13;
    adder_0_reduction_io_r_delay_15 <= adder_0_reduction_io_r_delay_14;
    adder_0_reduction_io_r_delay_16 <= adder_0_reduction_io_r_delay_15;
    adder_0_reduction_io_r_delay_17 <= adder_0_reduction_io_r_delay_16;
    adder_0_reduction_io_r_delay_18 <= adder_0_reduction_io_r_delay_17;
    adder_0_reduction_io_r_delay_19 <= adder_0_reduction_io_r_delay_18;
    adder_0_reduction_io_r_delay_20 <= adder_0_reduction_io_r_delay_19;
    adder_0_reduction_io_r_delay_21 <= adder_0_reduction_io_r_delay_20;
    adder_0_reduction_io_r_delay_22 <= adder_0_reduction_io_r_delay_21;
    adder_0_reduction_io_r_delay_23 <= adder_0_reduction_io_r_delay_22;
    adder_0_reduction_io_r_delay_24 <= adder_0_reduction_io_r_delay_23;
    adder_0_reduction_io_r_delay_25 <= adder_0_reduction_io_r_delay_24;
    adder_0_reduction_io_r_delay_26 <= adder_0_reduction_io_r_delay_25;
    adder_0_reduction_io_r_delay_27 <= adder_0_reduction_io_r_delay_26;
    adder_0_reduction_io_r_delay_28 <= adder_0_reduction_io_r_delay_27;
    adder_0_reduction_io_r_delay_29 <= adder_0_reduction_io_r_delay_28;
    adder_0_reduction_io_r_delay_30 <= adder_0_reduction_io_r_delay_29;
    adder_0_reduction_io_r_delay_31 <= adder_0_reduction_io_r_delay_30;
    adder_0_reduction_io_r_delay_32 <= adder_0_reduction_io_r_delay_31;
    adder_0_reduction_io_r_delay_33 <= adder_0_reduction_io_r_delay_32;
    adder_0_reduction_io_r_delay_34 <= adder_0_reduction_io_r_delay_33;
    adder_0_reduction_io_r_delay_35 <= adder_0_reduction_io_r_delay_34;
    adder_0_reduction_io_r_delay_36 <= adder_0_reduction_io_r_delay_35;
    adder_0_reduction_io_r_delay_37 <= adder_0_reduction_io_r_delay_36;
    adder_0_reduction_io_r_delay_38 <= adder_0_reduction_io_r_delay_37;
    adder_0_reduction_io_r_delay_39 <= adder_0_reduction_io_r_delay_38;
    adder_0_reduction_io_r_delay_40 <= adder_0_reduction_io_r_delay_39;
    adder_0_reduction_io_r_delay_41 <= adder_0_reduction_io_r_delay_40;
    adder_0_reduction_io_r_delay_42 <= adder_0_reduction_io_r_delay_41;
    adder_0_reduction_io_r_delay_43 <= adder_0_reduction_io_r_delay_42;
    adder_0_reduction_io_r_delay_44 <= adder_0_reduction_io_r_delay_43;
    adder_0_reduction_io_r_delay_45 <= adder_0_reduction_io_r_delay_44;
    adder_0_reduction_io_r_delay_46 <= adder_0_reduction_io_r_delay_45;
    adder_0_reduction_io_r_delay_47 <= adder_0_reduction_io_r_delay_46;
    adder_0_reduction_io_r_delay_48 <= adder_0_reduction_io_r_delay_47;
    adder_0_reduction_io_r_delay_49 <= adder_0_reduction_io_r_delay_48;
    adder_0_reduction_io_r_delay_50 <= adder_0_reduction_io_r_delay_49;
    adder_0_reduction_io_r_delay_51 <= adder_0_reduction_io_r_delay_50;
    adder_0_reduction_io_r_delay_52 <= adder_0_reduction_io_r_delay_51;
    adder_0_reduction_io_r_delay_53 <= adder_0_reduction_io_r_delay_52;
    adder_0_reduction_io_r_delay_54 <= adder_0_reduction_io_r_delay_53;
    adder_0_reduction_io_r_delay_55 <= adder_0_reduction_io_r_delay_54;
    adder_0_reduction_io_r_delay_56 <= adder_0_reduction_io_r_delay_55;
    adder_0_reduction_io_r_delay_57 <= adder_0_reduction_io_r_delay_56;
    adder_0_reduction_io_r_delay_58 <= adder_0_reduction_io_r_delay_57;
    adder_0_reduction_io_r_delay_59 <= adder_0_reduction_io_r_delay_58;
    adder_0_reduction_io_r_delay_60 <= adder_0_reduction_io_r_delay_59;
    adder_0_reduction_io_r_delay_61 <= adder_0_reduction_io_r_delay_60;
    adder_0_reduction_io_r_delay_62 <= adder_0_reduction_io_r_delay_61;
    adder_0_reduction_io_r_delay_63 <= adder_0_reduction_io_r_delay_62;
    adder_0_reduction_io_r_delay_64 <= adder_0_reduction_io_r_delay_63;
    adder_0_reduction_io_r_delay_65 <= adder_0_reduction_io_r_delay_64;
    adder_0_reduction_io_r_delay_66 <= adder_0_reduction_io_r_delay_65;
    adder_0_reduction_io_r_delay_67 <= adder_0_reduction_io_r_delay_66;
    adder_0_reduction_io_r_delay_68 <= adder_0_reduction_io_r_delay_67;
    adder_0_reduction_io_r_delay_69 <= adder_0_reduction_io_r_delay_68;
    adder_0_reduction_io_r_delay_70 <= adder_0_reduction_io_r_delay_69;
    adder_0_reduction_io_r_delay_71 <= adder_0_reduction_io_r_delay_70;
    adder_0_reduction_io_r_delay_72 <= adder_0_reduction_io_r_delay_71;
    adder_0_reduction_io_r_delay_73 <= adder_0_reduction_io_r_delay_72;
    adder_0_reduction_io_r_delay_74 <= adder_0_reduction_io_r_delay_73;
    adder_0_reduction_io_r_delay_75 <= adder_0_reduction_io_r_delay_74;
    adder_0_reduction_io_r_delay_76 <= adder_0_reduction_io_r_delay_75;
    R8 <= adder_0_reduction_io_r_delay_76;
    adder_0_sub_2_io_s_delay_1 <= sub_2_io_s;
    adder_0_sub_2_io_s_delay_2 <= adder_0_sub_2_io_s_delay_1;
    adder_0_sub_2_io_s_delay_3 <= adder_0_sub_2_io_s_delay_2;
    adder_0_sub_2_io_s_delay_4 <= adder_0_sub_2_io_s_delay_3;
    adder_0_sub_2_io_s_delay_5 <= adder_0_sub_2_io_s_delay_4;
    adder_0_sub_2_io_s_delay_6 <= adder_0_sub_2_io_s_delay_5;
    adder_0_sub_2_io_s_delay_7 <= adder_0_sub_2_io_s_delay_6;
    adder_0_sub_2_io_s_delay_8 <= adder_0_sub_2_io_s_delay_7;
    adder_0_sub_2_io_s_delay_9 <= adder_0_sub_2_io_s_delay_8;
    adder_0_sub_2_io_s_delay_10 <= adder_0_sub_2_io_s_delay_9;
    adder_0_sub_2_io_s_delay_11 <= adder_0_sub_2_io_s_delay_10;
    adder_0_sub_2_io_s_delay_12 <= adder_0_sub_2_io_s_delay_11;
    adder_0_sub_2_io_s_delay_13 <= adder_0_sub_2_io_s_delay_12;
    adder_0_sub_2_io_s_delay_14 <= adder_0_sub_2_io_s_delay_13;
    adder_0_sub_2_io_s_delay_15 <= adder_0_sub_2_io_s_delay_14;
    adder_0_sub_2_io_s_delay_16 <= adder_0_sub_2_io_s_delay_15;
    adder_0_sub_2_io_s_delay_17 <= adder_0_sub_2_io_s_delay_16;
    adder_0_sub_2_io_s_delay_18 <= adder_0_sub_2_io_s_delay_17;
    adder_0_sub_2_io_s_delay_19 <= adder_0_sub_2_io_s_delay_18;
    adder_0_sub_2_io_s_delay_20 <= adder_0_sub_2_io_s_delay_19;
    adder_0_sub_2_io_s_delay_21 <= adder_0_sub_2_io_s_delay_20;
    adder_0_sub_2_io_s_delay_22 <= adder_0_sub_2_io_s_delay_21;
    adder_0_sub_2_io_s_delay_23 <= adder_0_sub_2_io_s_delay_22;
    adder_0_sub_2_io_s_delay_24 <= adder_0_sub_2_io_s_delay_23;
    adder_0_sub_2_io_s_delay_25 <= adder_0_sub_2_io_s_delay_24;
    adder_0_sub_2_io_s_delay_26 <= adder_0_sub_2_io_s_delay_25;
    adder_0_sub_2_io_s_delay_27 <= adder_0_sub_2_io_s_delay_26;
    adder_0_sub_2_io_s_delay_28 <= adder_0_sub_2_io_s_delay_27;
    adder_0_sub_2_io_s_delay_29 <= adder_0_sub_2_io_s_delay_28;
    adder_0_sub_2_io_s_delay_30 <= adder_0_sub_2_io_s_delay_29;
    adder_0_sub_2_io_s_delay_31 <= adder_0_sub_2_io_s_delay_30;
    adder_0_sub_2_io_s_delay_32 <= adder_0_sub_2_io_s_delay_31;
    adder_0_sub_2_io_s_delay_33 <= adder_0_sub_2_io_s_delay_32;
    adder_0_sub_2_io_s_delay_34 <= adder_0_sub_2_io_s_delay_33;
    adder_0_sub_2_io_s_delay_35 <= adder_0_sub_2_io_s_delay_34;
    adder_0_sub_2_io_s_delay_36 <= adder_0_sub_2_io_s_delay_35;
    adder_0_sub_2_io_s_delay_37 <= adder_0_sub_2_io_s_delay_36;
    adder_0_sub_2_io_s_delay_38 <= adder_0_sub_2_io_s_delay_37;
    adder_0_sub_2_io_s_delay_39 <= adder_0_sub_2_io_s_delay_38;
    adder_0_sub_2_io_s_delay_40 <= adder_0_sub_2_io_s_delay_39;
    adder_0_sub_2_io_s_delay_41 <= adder_0_sub_2_io_s_delay_40;
    adder_0_sub_2_io_s_delay_42 <= adder_0_sub_2_io_s_delay_41;
    adder_0_sub_2_io_s_delay_43 <= adder_0_sub_2_io_s_delay_42;
    adder_0_sub_2_io_s_delay_44 <= adder_0_sub_2_io_s_delay_43;
    adder_0_sub_2_io_s_delay_45 <= adder_0_sub_2_io_s_delay_44;
    adder_0_sub_2_io_s_delay_46 <= adder_0_sub_2_io_s_delay_45;
    adder_0_sub_2_io_s_delay_47 <= adder_0_sub_2_io_s_delay_46;
    adder_0_sub_2_io_s_delay_48 <= adder_0_sub_2_io_s_delay_47;
    adder_0_sub_2_io_s_delay_49 <= adder_0_sub_2_io_s_delay_48;
    adder_0_sub_2_io_s_delay_50 <= adder_0_sub_2_io_s_delay_49;
    adder_0_sub_2_io_s_delay_51 <= adder_0_sub_2_io_s_delay_50;
    adder_0_sub_2_io_s_delay_52 <= adder_0_sub_2_io_s_delay_51;
    adder_0_sub_2_io_s_delay_53 <= adder_0_sub_2_io_s_delay_52;
    adder_0_sub_2_io_s_delay_54 <= adder_0_sub_2_io_s_delay_53;
    adder_0_sub_2_io_s_delay_55 <= adder_0_sub_2_io_s_delay_54;
    adder_0_sub_2_io_s_delay_56 <= adder_0_sub_2_io_s_delay_55;
    adder_0_sub_2_io_s_delay_57 <= adder_0_sub_2_io_s_delay_56;
    adder_0_sub_2_io_s_delay_58 <= adder_0_sub_2_io_s_delay_57;
    adder_0_sub_2_io_s_delay_59 <= adder_0_sub_2_io_s_delay_58;
    adder_0_sub_2_io_s_delay_60 <= adder_0_sub_2_io_s_delay_59;
    adder_0_sub_2_io_s_delay_61 <= adder_0_sub_2_io_s_delay_60;
    adder_0_sub_2_io_s_delay_62 <= adder_0_sub_2_io_s_delay_61;
    adder_0_sub_2_io_s_delay_63 <= adder_0_sub_2_io_s_delay_62;
    adder_0_sub_2_io_s_delay_64 <= adder_0_sub_2_io_s_delay_63;
    adder_0_sub_2_io_s_delay_65 <= adder_0_sub_2_io_s_delay_64;
    adder_0_sub_2_io_s_delay_66 <= adder_0_sub_2_io_s_delay_65;
    adder_0_sub_2_io_s_delay_67 <= adder_0_sub_2_io_s_delay_66;
    adder_0_sub_2_io_s_delay_68 <= adder_0_sub_2_io_s_delay_67;
    adder_0_sub_2_io_s_delay_69 <= adder_0_sub_2_io_s_delay_68;
    adder_0_sub_2_io_s_delay_70 <= adder_0_sub_2_io_s_delay_69;
    adder_0_sub_2_io_s_delay_71 <= adder_0_sub_2_io_s_delay_70;
    adder_0_sub_2_io_s_delay_72 <= adder_0_sub_2_io_s_delay_71;
    adder_0_sub_2_io_s_delay_73 <= adder_0_sub_2_io_s_delay_72;
    adder_0_sub_2_io_s_delay_74 <= adder_0_sub_2_io_s_delay_73;
    adder_0_sub_2_io_s_delay_75 <= adder_0_sub_2_io_s_delay_74;
    R9 <= adder_0_sub_2_io_s_delay_75;
    adder_0_add_3_io_s_delay_1 <= add_3_io_s;
    adder_0_add_3_io_s_delay_2 <= adder_0_add_3_io_s_delay_1;
    adder_0_add_3_io_s_delay_3 <= adder_0_add_3_io_s_delay_2;
    adder_0_add_3_io_s_delay_4 <= adder_0_add_3_io_s_delay_3;
    adder_0_add_3_io_s_delay_5 <= adder_0_add_3_io_s_delay_4;
    adder_0_add_3_io_s_delay_6 <= adder_0_add_3_io_s_delay_5;
    adder_0_add_3_io_s_delay_7 <= adder_0_add_3_io_s_delay_6;
    adder_0_add_3_io_s_delay_8 <= adder_0_add_3_io_s_delay_7;
    adder_0_add_3_io_s_delay_9 <= adder_0_add_3_io_s_delay_8;
    adder_0_add_3_io_s_delay_10 <= adder_0_add_3_io_s_delay_9;
    adder_0_add_3_io_s_delay_11 <= adder_0_add_3_io_s_delay_10;
    adder_0_add_3_io_s_delay_12 <= adder_0_add_3_io_s_delay_11;
    adder_0_add_3_io_s_delay_13 <= adder_0_add_3_io_s_delay_12;
    adder_0_add_3_io_s_delay_14 <= adder_0_add_3_io_s_delay_13;
    adder_0_add_3_io_s_delay_15 <= adder_0_add_3_io_s_delay_14;
    adder_0_add_3_io_s_delay_16 <= adder_0_add_3_io_s_delay_15;
    adder_0_add_3_io_s_delay_17 <= adder_0_add_3_io_s_delay_16;
    adder_0_add_3_io_s_delay_18 <= adder_0_add_3_io_s_delay_17;
    adder_0_add_3_io_s_delay_19 <= adder_0_add_3_io_s_delay_18;
    adder_0_add_3_io_s_delay_20 <= adder_0_add_3_io_s_delay_19;
    adder_0_add_3_io_s_delay_21 <= adder_0_add_3_io_s_delay_20;
    adder_0_add_3_io_s_delay_22 <= adder_0_add_3_io_s_delay_21;
    adder_0_add_3_io_s_delay_23 <= adder_0_add_3_io_s_delay_22;
    adder_0_add_3_io_s_delay_24 <= adder_0_add_3_io_s_delay_23;
    adder_0_add_3_io_s_delay_25 <= adder_0_add_3_io_s_delay_24;
    adder_0_add_3_io_s_delay_26 <= adder_0_add_3_io_s_delay_25;
    adder_0_add_3_io_s_delay_27 <= adder_0_add_3_io_s_delay_26;
    adder_0_add_3_io_s_delay_28 <= adder_0_add_3_io_s_delay_27;
    adder_0_add_3_io_s_delay_29 <= adder_0_add_3_io_s_delay_28;
    adder_0_add_3_io_s_delay_30 <= adder_0_add_3_io_s_delay_29;
    adder_0_add_3_io_s_delay_31 <= adder_0_add_3_io_s_delay_30;
    adder_0_add_3_io_s_delay_32 <= adder_0_add_3_io_s_delay_31;
    adder_0_add_3_io_s_delay_33 <= adder_0_add_3_io_s_delay_32;
    adder_0_add_3_io_s_delay_34 <= adder_0_add_3_io_s_delay_33;
    adder_0_add_3_io_s_delay_35 <= adder_0_add_3_io_s_delay_34;
    adder_0_add_3_io_s_delay_36 <= adder_0_add_3_io_s_delay_35;
    adder_0_add_3_io_s_delay_37 <= adder_0_add_3_io_s_delay_36;
    adder_0_add_3_io_s_delay_38 <= adder_0_add_3_io_s_delay_37;
    adder_0_add_3_io_s_delay_39 <= adder_0_add_3_io_s_delay_38;
    adder_0_add_3_io_s_delay_40 <= adder_0_add_3_io_s_delay_39;
    adder_0_add_3_io_s_delay_41 <= adder_0_add_3_io_s_delay_40;
    adder_0_add_3_io_s_delay_42 <= adder_0_add_3_io_s_delay_41;
    adder_0_add_3_io_s_delay_43 <= adder_0_add_3_io_s_delay_42;
    adder_0_add_3_io_s_delay_44 <= adder_0_add_3_io_s_delay_43;
    adder_0_add_3_io_s_delay_45 <= adder_0_add_3_io_s_delay_44;
    adder_0_add_3_io_s_delay_46 <= adder_0_add_3_io_s_delay_45;
    adder_0_add_3_io_s_delay_47 <= adder_0_add_3_io_s_delay_46;
    adder_0_add_3_io_s_delay_48 <= adder_0_add_3_io_s_delay_47;
    adder_0_add_3_io_s_delay_49 <= adder_0_add_3_io_s_delay_48;
    adder_0_add_3_io_s_delay_50 <= adder_0_add_3_io_s_delay_49;
    adder_0_add_3_io_s_delay_51 <= adder_0_add_3_io_s_delay_50;
    adder_0_add_3_io_s_delay_52 <= adder_0_add_3_io_s_delay_51;
    adder_0_add_3_io_s_delay_53 <= adder_0_add_3_io_s_delay_52;
    adder_0_add_3_io_s_delay_54 <= adder_0_add_3_io_s_delay_53;
    adder_0_add_3_io_s_delay_55 <= adder_0_add_3_io_s_delay_54;
    adder_0_add_3_io_s_delay_56 <= adder_0_add_3_io_s_delay_55;
    adder_0_add_3_io_s_delay_57 <= adder_0_add_3_io_s_delay_56;
    adder_0_add_3_io_s_delay_58 <= adder_0_add_3_io_s_delay_57;
    adder_0_add_3_io_s_delay_59 <= adder_0_add_3_io_s_delay_58;
    adder_0_add_3_io_s_delay_60 <= adder_0_add_3_io_s_delay_59;
    adder_0_add_3_io_s_delay_61 <= adder_0_add_3_io_s_delay_60;
    adder_0_add_3_io_s_delay_62 <= adder_0_add_3_io_s_delay_61;
    adder_0_add_3_io_s_delay_63 <= adder_0_add_3_io_s_delay_62;
    adder_0_add_3_io_s_delay_64 <= adder_0_add_3_io_s_delay_63;
    adder_0_add_3_io_s_delay_65 <= adder_0_add_3_io_s_delay_64;
    adder_0_add_3_io_s_delay_66 <= adder_0_add_3_io_s_delay_65;
    adder_0_add_3_io_s_delay_67 <= adder_0_add_3_io_s_delay_66;
    adder_0_add_3_io_s_delay_68 <= adder_0_add_3_io_s_delay_67;
    adder_0_add_3_io_s_delay_69 <= adder_0_add_3_io_s_delay_68;
    adder_0_add_3_io_s_delay_70 <= adder_0_add_3_io_s_delay_69;
    adder_0_add_3_io_s_delay_71 <= adder_0_add_3_io_s_delay_70;
    adder_0_add_3_io_s_delay_72 <= adder_0_add_3_io_s_delay_71;
    adder_0_add_3_io_s_delay_73 <= adder_0_add_3_io_s_delay_72;
    adder_0_add_3_io_s_delay_74 <= adder_0_add_3_io_s_delay_73;
    adder_0_add_3_io_s_delay_75 <= adder_0_add_3_io_s_delay_74;
    R12 <= adder_0_add_3_io_s_delay_75;
  end


endmodule

module DWSRFIFO (
  input               io_dataIn_0_valid,
  input      [376:0]  io_dataIn_0_payload_a_X,
  input      [376:0]  io_dataIn_0_payload_a_Y,
  input      [376:0]  io_dataIn_0_payload_a_Z,
  input      [376:0]  io_dataIn_0_payload_a_T,
  input      [376:0]  io_dataIn_0_payload_b_X,
  input      [376:0]  io_dataIn_0_payload_b_Y,
  input      [376:0]  io_dataIn_0_payload_b_Z,
  input      [376:0]  io_dataIn_0_payload_b_T,
  input      [16:0]   io_dataIn_0_payload_address,
  input               io_dataIn_1_valid,
  input      [376:0]  io_dataIn_1_payload_a_X,
  input      [376:0]  io_dataIn_1_payload_a_Y,
  input      [376:0]  io_dataIn_1_payload_a_Z,
  input      [376:0]  io_dataIn_1_payload_a_T,
  input      [376:0]  io_dataIn_1_payload_b_X,
  input      [376:0]  io_dataIn_1_payload_b_Y,
  input      [376:0]  io_dataIn_1_payload_b_Z,
  input      [376:0]  io_dataIn_1_payload_b_T,
  input      [16:0]   io_dataIn_1_payload_address,
  output              io_dataOut_valid,
  output     [376:0]  io_dataOut_payload_a_X,
  output     [376:0]  io_dataOut_payload_a_Y,
  output     [376:0]  io_dataOut_payload_a_Z,
  output     [376:0]  io_dataOut_payload_a_T,
  output     [376:0]  io_dataOut_payload_b_X,
  output     [376:0]  io_dataOut_payload_b_Y,
  output     [376:0]  io_dataOut_payload_b_Z,
  output     [376:0]  io_dataOut_payload_b_T,
  output     [16:0]   io_dataOut_payload_address,
  input               clk,
  input               resetn
);

  wire       [376:0]  ram_io_rData_a_X;
  wire       [376:0]  ram_io_rData_a_Y;
  wire       [376:0]  ram_io_rData_a_Z;
  wire       [376:0]  ram_io_rData_a_T;
  wire       [376:0]  ram_io_rData_b_X;
  wire       [376:0]  ram_io_rData_b_Y;
  wire       [376:0]  ram_io_rData_b_Z;
  wire       [376:0]  ram_io_rData_b_T;
  wire       [16:0]   ram_io_rData_address;
  wire       [7:0]    _zz_pushPtr_valueNext;
  wire       [0:0]    _zz_pushPtr_valueNext_1;
  wire       [7:0]    _zz_popPtr_valueNext;
  wire       [0:0]    _zz_popPtr_valueNext_1;
  reg                 pushPtr_willIncrement;
  wire                pushPtr_willClear;
  reg        [7:0]    pushPtr_valueNext;
  reg        [7:0]    pushPtr_value;
  reg                 pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  wire                popPtr_willClear;
  reg        [7:0]    popPtr_valueNext;
  reg        [7:0]    popPtr_value;
  reg                 popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  reg                 empty;
  reg                 _zz_io_dataOut_valid;
  reg                 _zz_io_dataOut_valid_1;
  reg                 _zz_io_dataOut_valid_2;
  reg                 _zz_io_dataOut_valid_3;
  reg                 io_dataIn_1_valid_delay_1;
  reg                 io_dataIn_1_valid_delay_2;
  reg                 io_dataIn_1_valid_delay_3;
  reg                 io_dataIn_1_valid_delay_4;
  reg        [376:0]  io_dataIn_1_payload_delay_1_a_X;
  reg        [376:0]  io_dataIn_1_payload_delay_1_a_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_1_a_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_1_a_T;
  reg        [376:0]  io_dataIn_1_payload_delay_1_b_X;
  reg        [376:0]  io_dataIn_1_payload_delay_1_b_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_1_b_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_1_b_T;
  reg        [16:0]   io_dataIn_1_payload_delay_1_address;
  reg        [376:0]  io_dataIn_1_payload_delay_2_a_X;
  reg        [376:0]  io_dataIn_1_payload_delay_2_a_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_2_a_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_2_a_T;
  reg        [376:0]  io_dataIn_1_payload_delay_2_b_X;
  reg        [376:0]  io_dataIn_1_payload_delay_2_b_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_2_b_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_2_b_T;
  reg        [16:0]   io_dataIn_1_payload_delay_2_address;
  reg        [376:0]  io_dataIn_1_payload_delay_3_a_X;
  reg        [376:0]  io_dataIn_1_payload_delay_3_a_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_3_a_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_3_a_T;
  reg        [376:0]  io_dataIn_1_payload_delay_3_b_X;
  reg        [376:0]  io_dataIn_1_payload_delay_3_b_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_3_b_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_3_b_T;
  reg        [16:0]   io_dataIn_1_payload_delay_3_address;
  reg        [376:0]  io_dataIn_1_payload_delay_4_a_X;
  reg        [376:0]  io_dataIn_1_payload_delay_4_a_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_4_a_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_4_a_T;
  reg        [376:0]  io_dataIn_1_payload_delay_4_b_X;
  reg        [376:0]  io_dataIn_1_payload_delay_4_b_Y;
  reg        [376:0]  io_dataIn_1_payload_delay_4_b_Z;
  reg        [376:0]  io_dataIn_1_payload_delay_4_b_T;
  reg        [16:0]   io_dataIn_1_payload_delay_4_address;
  wire                when_DWSRFIFO_l41;

  assign _zz_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign _zz_pushPtr_valueNext = {7'd0, _zz_pushPtr_valueNext_1};
  assign _zz_popPtr_valueNext_1 = popPtr_willIncrement;
  assign _zz_popPtr_valueNext = {7'd0, _zz_popPtr_valueNext_1};
  SDPRAM ram (
    .io_we            (io_dataIn_0_valid                ), //i
    .io_wAddress      (pushPtr_value[7:0]               ), //i
    .io_wData_a_X     (io_dataIn_0_payload_a_X[376:0]   ), //i
    .io_wData_a_Y     (io_dataIn_0_payload_a_Y[376:0]   ), //i
    .io_wData_a_Z     (io_dataIn_0_payload_a_Z[376:0]   ), //i
    .io_wData_a_T     (io_dataIn_0_payload_a_T[376:0]   ), //i
    .io_wData_b_X     (io_dataIn_0_payload_b_X[376:0]   ), //i
    .io_wData_b_Y     (io_dataIn_0_payload_b_Y[376:0]   ), //i
    .io_wData_b_Z     (io_dataIn_0_payload_b_Z[376:0]   ), //i
    .io_wData_b_T     (io_dataIn_0_payload_b_T[376:0]   ), //i
    .io_wData_address (io_dataIn_0_payload_address[16:0]), //i
    .io_re            (1'b1                             ), //i
    .io_rAddress      (popPtr_value[7:0]                ), //i
    .io_rData_a_X     (ram_io_rData_a_X[376:0]          ), //o
    .io_rData_a_Y     (ram_io_rData_a_Y[376:0]          ), //o
    .io_rData_a_Z     (ram_io_rData_a_Z[376:0]          ), //o
    .io_rData_a_T     (ram_io_rData_a_T[376:0]          ), //o
    .io_rData_b_X     (ram_io_rData_b_X[376:0]          ), //o
    .io_rData_b_Y     (ram_io_rData_b_Y[376:0]          ), //o
    .io_rData_b_Z     (ram_io_rData_b_Z[376:0]          ), //o
    .io_rData_b_T     (ram_io_rData_b_T[376:0]          ), //o
    .io_rData_address (ram_io_rData_address[16:0]       ), //o
    .clk              (clk                              ), //i
    .resetn           (resetn                           )  //i
  );
  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(io_dataIn_0_valid) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  assign pushPtr_willClear = 1'b0;
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    pushPtr_valueNext = (pushPtr_value + _zz_pushPtr_valueNext);
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 8'h0;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(when_DWSRFIFO_l41) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  assign popPtr_willClear = 1'b0;
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    popPtr_valueNext = (popPtr_value + _zz_popPtr_valueNext);
    if(popPtr_willClear) begin
      popPtr_valueNext = 8'h0;
    end
  end

  assign io_dataOut_valid = _zz_io_dataOut_valid_3;
  assign io_dataOut_payload_a_X = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_a_X : ram_io_rData_a_X);
  assign io_dataOut_payload_a_Y = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_a_Y : ram_io_rData_a_Y);
  assign io_dataOut_payload_a_Z = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_a_Z : ram_io_rData_a_Z);
  assign io_dataOut_payload_a_T = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_a_T : ram_io_rData_a_T);
  assign io_dataOut_payload_b_X = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_b_X : ram_io_rData_b_X);
  assign io_dataOut_payload_b_Y = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_b_Y : ram_io_rData_b_Y);
  assign io_dataOut_payload_b_Z = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_b_Z : ram_io_rData_b_Z);
  assign io_dataOut_payload_b_T = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_b_T : ram_io_rData_b_T);
  assign io_dataOut_payload_address = (io_dataIn_1_valid_delay_4 ? io_dataIn_1_payload_delay_4_address : ram_io_rData_address);
  assign when_DWSRFIFO_l41 = ((! empty) && (! io_dataIn_1_valid));
  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      pushPtr_value <= 8'h0;
      pushPtr_willOverflowIfInc <= 1'b0;
      popPtr_value <= 8'h0;
      popPtr_willOverflowIfInc <= 1'b0;
      empty <= 1'b1;
      _zz_io_dataOut_valid <= 1'b0;
      _zz_io_dataOut_valid_1 <= 1'b0;
      _zz_io_dataOut_valid_2 <= 1'b0;
      _zz_io_dataOut_valid_3 <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      pushPtr_willOverflowIfInc <= (pushPtr_valueNext == 8'hff);
      popPtr_value <= popPtr_valueNext;
      popPtr_willOverflowIfInc <= (popPtr_valueNext == 8'hff);
      empty <= (pushPtr_value == popPtr_valueNext);
      _zz_io_dataOut_valid <= ((! empty) || io_dataIn_1_valid);
      _zz_io_dataOut_valid_1 <= _zz_io_dataOut_valid;
      _zz_io_dataOut_valid_2 <= _zz_io_dataOut_valid_1;
      _zz_io_dataOut_valid_3 <= _zz_io_dataOut_valid_2;
    end
  end

  always @(posedge clk) begin
    io_dataIn_1_valid_delay_1 <= io_dataIn_1_valid;
    io_dataIn_1_valid_delay_2 <= io_dataIn_1_valid_delay_1;
    io_dataIn_1_valid_delay_3 <= io_dataIn_1_valid_delay_2;
    io_dataIn_1_valid_delay_4 <= io_dataIn_1_valid_delay_3;
    io_dataIn_1_payload_delay_1_a_X <= io_dataIn_1_payload_a_X;
    io_dataIn_1_payload_delay_1_a_Y <= io_dataIn_1_payload_a_Y;
    io_dataIn_1_payload_delay_1_a_Z <= io_dataIn_1_payload_a_Z;
    io_dataIn_1_payload_delay_1_a_T <= io_dataIn_1_payload_a_T;
    io_dataIn_1_payload_delay_1_b_X <= io_dataIn_1_payload_b_X;
    io_dataIn_1_payload_delay_1_b_Y <= io_dataIn_1_payload_b_Y;
    io_dataIn_1_payload_delay_1_b_Z <= io_dataIn_1_payload_b_Z;
    io_dataIn_1_payload_delay_1_b_T <= io_dataIn_1_payload_b_T;
    io_dataIn_1_payload_delay_1_address <= io_dataIn_1_payload_address;
    io_dataIn_1_payload_delay_2_a_X <= io_dataIn_1_payload_delay_1_a_X;
    io_dataIn_1_payload_delay_2_a_Y <= io_dataIn_1_payload_delay_1_a_Y;
    io_dataIn_1_payload_delay_2_a_Z <= io_dataIn_1_payload_delay_1_a_Z;
    io_dataIn_1_payload_delay_2_a_T <= io_dataIn_1_payload_delay_1_a_T;
    io_dataIn_1_payload_delay_2_b_X <= io_dataIn_1_payload_delay_1_b_X;
    io_dataIn_1_payload_delay_2_b_Y <= io_dataIn_1_payload_delay_1_b_Y;
    io_dataIn_1_payload_delay_2_b_Z <= io_dataIn_1_payload_delay_1_b_Z;
    io_dataIn_1_payload_delay_2_b_T <= io_dataIn_1_payload_delay_1_b_T;
    io_dataIn_1_payload_delay_2_address <= io_dataIn_1_payload_delay_1_address;
    io_dataIn_1_payload_delay_3_a_X <= io_dataIn_1_payload_delay_2_a_X;
    io_dataIn_1_payload_delay_3_a_Y <= io_dataIn_1_payload_delay_2_a_Y;
    io_dataIn_1_payload_delay_3_a_Z <= io_dataIn_1_payload_delay_2_a_Z;
    io_dataIn_1_payload_delay_3_a_T <= io_dataIn_1_payload_delay_2_a_T;
    io_dataIn_1_payload_delay_3_b_X <= io_dataIn_1_payload_delay_2_b_X;
    io_dataIn_1_payload_delay_3_b_Y <= io_dataIn_1_payload_delay_2_b_Y;
    io_dataIn_1_payload_delay_3_b_Z <= io_dataIn_1_payload_delay_2_b_Z;
    io_dataIn_1_payload_delay_3_b_T <= io_dataIn_1_payload_delay_2_b_T;
    io_dataIn_1_payload_delay_3_address <= io_dataIn_1_payload_delay_2_address;
    io_dataIn_1_payload_delay_4_a_X <= io_dataIn_1_payload_delay_3_a_X;
    io_dataIn_1_payload_delay_4_a_Y <= io_dataIn_1_payload_delay_3_a_Y;
    io_dataIn_1_payload_delay_4_a_Z <= io_dataIn_1_payload_delay_3_a_Z;
    io_dataIn_1_payload_delay_4_a_T <= io_dataIn_1_payload_delay_3_a_T;
    io_dataIn_1_payload_delay_4_b_X <= io_dataIn_1_payload_delay_3_b_X;
    io_dataIn_1_payload_delay_4_b_Y <= io_dataIn_1_payload_delay_3_b_Y;
    io_dataIn_1_payload_delay_4_b_Z <= io_dataIn_1_payload_delay_3_b_Z;
    io_dataIn_1_payload_delay_4_b_T <= io_dataIn_1_payload_delay_3_b_T;
    io_dataIn_1_payload_delay_4_address <= io_dataIn_1_payload_delay_3_address;
  end


endmodule

module DataRam (
  input               io_we_0,
  input               io_we_1,
  input      [16:0]   io_address_0,
  input      [16:0]   io_address_1,
  input      [376:0]  io_wData_0_X,
  input      [376:0]  io_wData_0_Y,
  input      [376:0]  io_wData_0_Z,
  input      [376:0]  io_wData_0_T,
  input      [376:0]  io_wData_1_X,
  input      [376:0]  io_wData_1_Y,
  input      [376:0]  io_wData_1_Z,
  input      [376:0]  io_wData_1_T,
  input               io_state_0,
  input               io_state_1,
  output     [376:0]  io_rData_0_X,
  output     [376:0]  io_rData_0_Y,
  output     [376:0]  io_rData_0_Z,
  output     [376:0]  io_rData_0_T,
  output     [376:0]  io_rData_1_X,
  output     [376:0]  io_rData_1_Y,
  output     [376:0]  io_rData_1_Z,
  output     [376:0]  io_rData_1_T,
  input      [376:0]  io_pInit_X,
  input      [376:0]  io_pInit_Y,
  input      [376:0]  io_pInit_Z,
  input      [376:0]  io_pInit_T,
  input               clk,
  input               resetn
);

  wire       [376:0]  ram_io_rData_0_X;
  wire       [376:0]  ram_io_rData_0_Y;
  wire       [376:0]  ram_io_rData_0_Z;
  wire       [376:0]  ram_io_rData_0_T;
  wire       [376:0]  ram_io_rData_1_X;
  wire       [376:0]  ram_io_rData_1_Y;
  wire       [376:0]  ram_io_rData_1_Z;
  wire       [376:0]  ram_io_rData_1_T;
  reg        [376:0]  _zz_io_rData_0_X;
  reg        [376:0]  _zz_io_rData_0_Y;
  reg        [376:0]  _zz_io_rData_0_Z;
  reg        [376:0]  _zz_io_rData_0_T;
  reg        [376:0]  _zz_io_rData_1_X;
  reg        [376:0]  _zz_io_rData_1_Y;
  reg        [376:0]  _zz_io_rData_1_Z;
  reg        [376:0]  _zz_io_rData_1_T;

  TDPRAM ram (
    .io_we_0      (io_we_0                ), //i
    .io_we_1      (io_we_1                ), //i
    .io_address_0 (io_address_0[16:0]     ), //i
    .io_address_1 (io_address_1[16:0]     ), //i
    .io_wData_0_X (io_wData_0_X[376:0]    ), //i
    .io_wData_0_Y (io_wData_0_Y[376:0]    ), //i
    .io_wData_0_Z (io_wData_0_Z[376:0]    ), //i
    .io_wData_0_T (io_wData_0_T[376:0]    ), //i
    .io_wData_1_X (io_wData_1_X[376:0]    ), //i
    .io_wData_1_Y (io_wData_1_Y[376:0]    ), //i
    .io_wData_1_Z (io_wData_1_Z[376:0]    ), //i
    .io_wData_1_T (io_wData_1_T[376:0]    ), //i
    .io_ce_0      (1'b1                   ), //i
    .io_ce_1      (1'b1                   ), //i
    .io_rData_0_X (ram_io_rData_0_X[376:0]), //o
    .io_rData_0_Y (ram_io_rData_0_Y[376:0]), //o
    .io_rData_0_Z (ram_io_rData_0_Z[376:0]), //o
    .io_rData_0_T (ram_io_rData_0_T[376:0]), //o
    .io_rData_1_X (ram_io_rData_1_X[376:0]), //o
    .io_rData_1_Y (ram_io_rData_1_Y[376:0]), //o
    .io_rData_1_Z (ram_io_rData_1_Z[376:0]), //o
    .io_rData_1_T (ram_io_rData_1_T[376:0]), //o
    .clk          (clk                    ), //i
    .resetn       (resetn                 )  //i
  );
  assign io_rData_0_X = _zz_io_rData_0_X;
  assign io_rData_0_Y = _zz_io_rData_0_Y;
  assign io_rData_0_Z = _zz_io_rData_0_Z;
  assign io_rData_0_T = _zz_io_rData_0_T;
  assign io_rData_1_X = _zz_io_rData_1_X;
  assign io_rData_1_Y = _zz_io_rData_1_Y;
  assign io_rData_1_Z = _zz_io_rData_1_Z;
  assign io_rData_1_T = _zz_io_rData_1_T;
  always @(posedge clk) begin
    _zz_io_rData_0_X <= (io_state_0 ? ram_io_rData_0_X : io_pInit_X);
    _zz_io_rData_0_Y <= (io_state_0 ? ram_io_rData_0_Y : io_pInit_Y);
    _zz_io_rData_0_Z <= (io_state_0 ? ram_io_rData_0_Z : io_pInit_Z);
    _zz_io_rData_0_T <= (io_state_0 ? ram_io_rData_0_T : io_pInit_T);
    _zz_io_rData_1_X <= (io_state_1 ? ram_io_rData_1_X : io_pInit_X);
    _zz_io_rData_1_Y <= (io_state_1 ? ram_io_rData_1_Y : io_pInit_Y);
    _zz_io_rData_1_Z <= (io_state_1 ? ram_io_rData_1_Z : io_pInit_Z);
    _zz_io_rData_1_T <= (io_state_1 ? ram_io_rData_1_T : io_pInit_T);
  end


endmodule

module StateRam (
  input               io_we_0,
  input               io_we_1,
  input      [16:0]   io_address_0,
  input      [16:0]   io_address_1,
  output              io_state_0,
  output              io_state_1,
  input               io_flush,
  input      [16:0]   io_flushCnt,
  input               clk,
  input               resetn
);

  reg                 rams_0_0_io_we;
  reg        [16:0]   rams_0_0_io_wAddress;
  reg                 rams_0_0_io_wData;
  reg                 rams_0_1_io_we;
  reg        [16:0]   rams_0_1_io_wAddress;
  reg                 rams_0_1_io_wData;
  reg                 rams_1_0_io_we;
  reg        [16:0]   rams_1_0_io_wAddress;
  reg                 rams_1_0_io_wData;
  reg                 rams_1_1_io_we;
  reg        [16:0]   rams_1_1_io_wAddress;
  reg                 rams_1_1_io_wData;
  wire                rams_0_0_io_rData;
  wire                rams_0_1_io_rData;
  wire                rams_1_0_io_rData;
  wire                rams_1_1_io_rData;
  reg                 io_we_delay_1_0;
  reg                 io_we_delay_1_1;
  reg                 io_we_delay_2_0;
  reg                 io_we_delay_2_1;
  reg                 io_we_delay_3_0;
  reg                 io_we_delay_3_1;
  reg                 readArea_we_0;
  reg                 readArea_we_1;
  reg        [16:0]   io_address_regNext_0;
  reg        [16:0]   io_address_regNext_1;
  wire       [16:0]   readArea_address_0_0;
  wire       [16:0]   readArea_address_0_1;
  reg        [16:0]   readArea_address_1_0;
  reg        [16:0]   readArea_address_1_1;
  reg        [16:0]   readArea_address_2_0;
  reg        [16:0]   readArea_address_2_1;
  reg        [16:0]   readArea_address_3_0;
  reg        [16:0]   readArea_address_3_1;
  reg                 readArea_needFlip_0_0_0;
  reg                 readArea_needFlip_0_0_1;
  reg                 readArea_needFlip_0_1_0;
  reg                 readArea_needFlip_0_1_1;
  reg                 readArea_needFlip_1_0_0;
  reg                 readArea_needFlip_1_0_1;
  reg                 readArea_needFlip_1_1_0;
  reg                 readArea_needFlip_1_1_1;
  reg                 readArea_needFlip_2_0_0;
  reg                 readArea_needFlip_2_0_1;
  reg                 readArea_needFlip_2_1_0;
  reg                 readArea_needFlip_2_1_1;
  reg        [16:0]   io_address_0_regNext;
  reg        [16:0]   io_address_0_regNext_1;
  reg        [16:0]   io_address_1_regNext;
  reg        [16:0]   io_address_1_regNext_1;
  reg                 _zz_io_state_0;
  reg                 _zz_io_state_1;
  reg                 io_flush_regNext;
  reg        [16:0]   io_flushCnt_regNext;
  reg        [16:0]   io_flushCnt_regNext_1;
  reg        [16:0]   io_flushCnt_regNext_2;
  reg        [16:0]   io_flushCnt_regNext_3;

  SDPRAM_1 rams_0_0 (
    .io_we       (rams_0_0_io_we            ), //i
    .io_wAddress (rams_0_0_io_wAddress[16:0]), //i
    .io_wData    (rams_0_0_io_wData         ), //i
    .io_re       (1'b1                      ), //i
    .io_rAddress (io_address_0_regNext[16:0]), //i
    .io_rData    (rams_0_0_io_rData         ), //o
    .clk         (clk                       ), //i
    .resetn      (resetn                    )  //i
  );
  SDPRAM_1 rams_0_1 (
    .io_we       (rams_0_1_io_we            ), //i
    .io_wAddress (rams_0_1_io_wAddress[16:0]), //i
    .io_wData    (rams_0_1_io_wData         ), //i
    .io_re       (1'b1                      ), //i
    .io_rAddress (io_address_1_regNext[16:0]), //i
    .io_rData    (rams_0_1_io_rData         ), //o
    .clk         (clk                       ), //i
    .resetn      (resetn                    )  //i
  );
  SDPRAM_1 rams_1_0 (
    .io_we       (rams_1_0_io_we              ), //i
    .io_wAddress (rams_1_0_io_wAddress[16:0]  ), //i
    .io_wData    (rams_1_0_io_wData           ), //i
    .io_re       (1'b1                        ), //i
    .io_rAddress (io_address_0_regNext_1[16:0]), //i
    .io_rData    (rams_1_0_io_rData           ), //o
    .clk         (clk                         ), //i
    .resetn      (resetn                      )  //i
  );
  SDPRAM_1 rams_1_1 (
    .io_we       (rams_1_1_io_we              ), //i
    .io_wAddress (rams_1_1_io_wAddress[16:0]  ), //i
    .io_wData    (rams_1_1_io_wData           ), //i
    .io_re       (1'b1                        ), //i
    .io_rAddress (io_address_1_regNext_1[16:0]), //i
    .io_rData    (rams_1_1_io_rData           ), //o
    .clk         (clk                         ), //i
    .resetn      (resetn                      )  //i
  );
  assign readArea_address_0_0 = io_address_regNext_0;
  assign readArea_address_0_1 = io_address_regNext_1;
  assign io_state_0 = _zz_io_state_0;
  assign io_state_1 = _zz_io_state_1;
  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_0_io_wAddress = io_flushCnt_regNext;
    end else begin
      rams_0_0_io_wAddress = readArea_address_3_0;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_1_io_wAddress = io_flushCnt_regNext_1;
    end else begin
      rams_0_1_io_wAddress = readArea_address_3_0;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_0_io_wAddress = io_flushCnt_regNext_2;
    end else begin
      rams_1_0_io_wAddress = readArea_address_3_1;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_1_io_wAddress = io_flushCnt_regNext_3;
    end else begin
      rams_1_1_io_wAddress = readArea_address_3_1;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_0_io_wData = 1'b0;
    end else begin
      rams_0_0_io_wData = (! (rams_0_0_io_rData ^ readArea_needFlip_2_0_0));
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_1_io_wData = 1'b0;
    end else begin
      rams_0_1_io_wData = (! (rams_0_0_io_rData ^ readArea_needFlip_2_0_0));
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_0_io_wData = 1'b0;
    end else begin
      rams_1_0_io_wData = (! (rams_1_1_io_rData ^ readArea_needFlip_2_1_1));
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_1_io_wData = 1'b0;
    end else begin
      rams_1_1_io_wData = (! (rams_1_1_io_rData ^ readArea_needFlip_2_1_1));
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_0_io_we = 1'b1;
    end else begin
      rams_0_0_io_we = readArea_we_0;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_0_1_io_we = 1'b1;
    end else begin
      rams_0_1_io_we = readArea_we_0;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_0_io_we = 1'b1;
    end else begin
      rams_1_0_io_we = readArea_we_1;
    end
  end

  always @(*) begin
    if(io_flush_regNext) begin
      rams_1_1_io_we = 1'b1;
    end else begin
      rams_1_1_io_we = readArea_we_1;
    end
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      io_we_delay_1_0 <= 1'b0;
      io_we_delay_1_1 <= 1'b0;
      io_we_delay_2_0 <= 1'b0;
      io_we_delay_2_1 <= 1'b0;
      io_we_delay_3_0 <= 1'b0;
      io_we_delay_3_1 <= 1'b0;
      readArea_we_0 <= 1'b0;
      readArea_we_1 <= 1'b0;
    end else begin
      io_we_delay_1_0 <= io_we_0;
      io_we_delay_1_1 <= io_we_1;
      io_we_delay_2_0 <= io_we_delay_1_0;
      io_we_delay_2_1 <= io_we_delay_1_1;
      io_we_delay_3_0 <= io_we_delay_2_0;
      io_we_delay_3_1 <= io_we_delay_2_1;
      readArea_we_0 <= io_we_delay_3_0;
      readArea_we_1 <= io_we_delay_3_1;
    end
  end

  always @(posedge clk) begin
    io_address_regNext_0 <= io_address_0;
    io_address_regNext_1 <= io_address_1;
    readArea_address_1_0 <= readArea_address_0_0;
    readArea_address_1_1 <= readArea_address_0_1;
    readArea_address_2_0 <= readArea_address_1_0;
    readArea_address_2_1 <= readArea_address_1_1;
    readArea_address_3_0 <= readArea_address_2_0;
    readArea_address_3_1 <= readArea_address_2_1;
    io_address_0_regNext <= io_address_0;
    io_address_0_regNext_1 <= io_address_0;
    io_address_1_regNext <= io_address_1;
    io_address_1_regNext_1 <= io_address_1;
    readArea_needFlip_0_0_0 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_0_0)) ^ 1'b0);
    readArea_needFlip_0_0_1 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_0_1)) ^ 1'b0);
    readArea_needFlip_0_1_0 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_0_0)) ^ 1'b0);
    readArea_needFlip_0_1_1 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_0_1)) ^ 1'b0);
    readArea_needFlip_1_0_0 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_1_0)) ^ readArea_needFlip_0_0_0);
    readArea_needFlip_1_0_1 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_1_1)) ^ readArea_needFlip_0_0_1);
    readArea_needFlip_1_1_0 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_1_0)) ^ readArea_needFlip_0_1_0);
    readArea_needFlip_1_1_1 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_1_1)) ^ readArea_needFlip_0_1_1);
    readArea_needFlip_2_0_0 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_2_0)) ^ readArea_needFlip_1_0_0);
    readArea_needFlip_2_0_1 <= ((readArea_we_0 && (readArea_address_3_0 == readArea_address_2_1)) ^ readArea_needFlip_1_0_1);
    readArea_needFlip_2_1_0 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_2_0)) ^ readArea_needFlip_1_1_0);
    readArea_needFlip_2_1_1 <= ((readArea_we_1 && (readArea_address_3_1 == readArea_address_2_1)) ^ readArea_needFlip_1_1_1);
    _zz_io_state_0 <= ((rams_0_0_io_rData ^ rams_1_0_io_rData) ^ (readArea_needFlip_2_0_0 ^ readArea_needFlip_2_1_0));
    _zz_io_state_1 <= ((rams_0_1_io_rData ^ rams_1_1_io_rData) ^ (readArea_needFlip_2_0_1 ^ readArea_needFlip_2_1_1));
    io_flush_regNext <= io_flush;
  end

  always @(posedge clk) begin
    io_flushCnt_regNext <= io_flushCnt;
    io_flushCnt_regNext_1 <= io_flushCnt;
    io_flushCnt_regNext_2 <= io_flushCnt;
    io_flushCnt_regNext_3 <= io_flushCnt;
  end


endmodule

module BADD (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  input               io_c,
  output reg [377:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [376:0]  _zz__zz_io_s_1;
  wire       [64:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [376:0]  _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_10;
  wire       [64:0]   _zz__zz_io_s_10_1;
  wire       [0:0]    _zz__zz_io_s_10_2;
  wire       [376:0]  _zz__zz_io_s_19;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [376:0]  _zz__zz_io_s_30;
  wire       [64:0]   _zz__zz_io_s_33;
  wire       [64:0]   _zz__zz_io_s_33_1;
  wire       [0:0]    _zz__zz_io_s_33_2;
  wire       [376:0]  _zz__zz_io_s_42;
  wire       [64:0]   _zz__zz_io_s_46;
  wire       [64:0]   _zz__zz_io_s_46_1;
  wire       [0:0]    _zz__zz_io_s_46_2;
  wire       [376:0]  _zz__zz_io_s_55;
  wire       [57:0]   _zz__zz_io_s_60;
  wire       [57:0]   _zz__zz_io_s_60_1;
  wire       [0:0]    _zz__zz_io_s_60_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  wire       [64:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg                 _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg        [63:0]   _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg        [63:0]   _zz_io_s_25;
  reg                 _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg        [63:0]   _zz_io_s_29;
  reg        [63:0]   _zz_io_s_30;
  reg        [63:0]   _zz_io_s_31;
  reg        [63:0]   _zz_io_s_32;
  wire       [64:0]   _zz_io_s_33;
  reg        [63:0]   _zz_io_s_34;
  reg        [63:0]   _zz_io_s_35;
  reg        [63:0]   _zz_io_s_36;
  reg                 _zz_io_s_37;
  reg        [63:0]   _zz_io_s_38;
  reg        [63:0]   _zz_io_s_39;
  reg        [63:0]   _zz_io_s_40;
  reg        [63:0]   _zz_io_s_41;
  reg        [63:0]   _zz_io_s_42;
  reg        [63:0]   _zz_io_s_43;
  reg        [63:0]   _zz_io_s_44;
  reg        [63:0]   _zz_io_s_45;
  wire       [64:0]   _zz_io_s_46;
  reg        [63:0]   _zz_io_s_47;
  reg        [63:0]   _zz_io_s_48;
  reg                 _zz_io_s_49;
  reg        [56:0]   _zz_io_s_50;
  reg        [56:0]   _zz_io_s_51;
  reg        [56:0]   _zz_io_s_52;
  reg        [56:0]   _zz_io_s_53;
  reg        [56:0]   _zz_io_s_54;
  reg        [56:0]   _zz_io_s_55;
  reg        [56:0]   _zz_io_s_56;
  reg        [56:0]   _zz_io_s_57;
  reg        [56:0]   _zz_io_s_58;
  reg        [56:0]   _zz_io_s_59;
  wire       [57:0]   _zz_io_s_60;
  reg        [56:0]   _zz_io_s_61;
  reg                 _zz_io_s_62;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,_zz__zz_io_s_1[63 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {64'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_9 = (~ io_b);
  assign _zz__zz_io_s_10 = ({1'b0,_zz_io_s_8} + {1'b0,_zz_io_s_9});
  assign _zz__zz_io_s_10_2 = _zz_io_s_7;
  assign _zz__zz_io_s_10_1 = {64'd0, _zz__zz_io_s_10_2};
  assign _zz__zz_io_s_19 = (~ io_b);
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_18} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_16;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_30 = (~ io_b);
  assign _zz__zz_io_s_33 = ({1'b0,_zz_io_s_29} + {1'b0,_zz_io_s_32});
  assign _zz__zz_io_s_33_2 = _zz_io_s_26;
  assign _zz__zz_io_s_33_1 = {64'd0, _zz__zz_io_s_33_2};
  assign _zz__zz_io_s_42 = (~ io_b);
  assign _zz__zz_io_s_46 = ({1'b0,_zz_io_s_41} + {1'b0,_zz_io_s_45});
  assign _zz__zz_io_s_46_2 = _zz_io_s_37;
  assign _zz__zz_io_s_46_1 = {64'd0, _zz__zz_io_s_46_2};
  assign _zz__zz_io_s_55 = (~ io_b);
  assign _zz__zz_io_s_60 = ({1'b0,_zz_io_s_54} + {1'b0,_zz_io_s_59});
  assign _zz__zz_io_s_60_2 = _zz_io_s_49;
  assign _zz__zz_io_s_60_1 = {57'd0, _zz__zz_io_s_60_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_6;
    io_s[127 : 64] = _zz_io_s_15;
    io_s[191 : 128] = _zz_io_s_25;
    io_s[255 : 192] = _zz_io_s_36;
    io_s[319 : 256] = _zz_io_s_48;
    io_s[376 : 320] = _zz_io_s_61;
    io_s[377] = (! _zz_io_s_62);
  end

  assign _zz_io_s_10 = (_zz__zz_io_s_10 + _zz__zz_io_s_10_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_33 = (_zz__zz_io_s_33 + _zz__zz_io_s_33_1);
  assign _zz_io_s_46 = (_zz__zz_io_s_46 + _zz__zz_io_s_46_1);
  assign _zz_io_s_60 = (_zz__zz_io_s_60 + _zz__zz_io_s_60_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= _zz_io_s[64];
    _zz_io_s_8 <= io_a[127 : 64];
    _zz_io_s_9 <= _zz__zz_io_s_9[127 : 64];
    _zz_io_s_11 <= _zz_io_s_10[63:0];
    _zz_io_s_12 <= _zz_io_s_11;
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= _zz_io_s_10[64];
    _zz_io_s_17 <= io_a[191 : 128];
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= _zz__zz_io_s_19[191 : 128];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_22;
    _zz_io_s_24 <= _zz_io_s_23;
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_21[64];
    _zz_io_s_27 <= io_a[255 : 192];
    _zz_io_s_28 <= _zz_io_s_27;
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz__zz_io_s_30[255 : 192];
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_32 <= _zz_io_s_31;
    _zz_io_s_34 <= _zz_io_s_33[63:0];
    _zz_io_s_35 <= _zz_io_s_34;
    _zz_io_s_36 <= _zz_io_s_35;
    _zz_io_s_37 <= _zz_io_s_33[64];
    _zz_io_s_38 <= io_a[319 : 256];
    _zz_io_s_39 <= _zz_io_s_38;
    _zz_io_s_40 <= _zz_io_s_39;
    _zz_io_s_41 <= _zz_io_s_40;
    _zz_io_s_42 <= _zz__zz_io_s_42[319 : 256];
    _zz_io_s_43 <= _zz_io_s_42;
    _zz_io_s_44 <= _zz_io_s_43;
    _zz_io_s_45 <= _zz_io_s_44;
    _zz_io_s_47 <= _zz_io_s_46[63:0];
    _zz_io_s_48 <= _zz_io_s_47;
    _zz_io_s_49 <= _zz_io_s_46[64];
    _zz_io_s_50 <= io_a[376 : 320];
    _zz_io_s_51 <= _zz_io_s_50;
    _zz_io_s_52 <= _zz_io_s_51;
    _zz_io_s_53 <= _zz_io_s_52;
    _zz_io_s_54 <= _zz_io_s_53;
    _zz_io_s_55 <= _zz__zz_io_s_55[376 : 320];
    _zz_io_s_56 <= _zz_io_s_55;
    _zz_io_s_57 <= _zz_io_s_56;
    _zz_io_s_58 <= _zz_io_s_57;
    _zz_io_s_59 <= _zz_io_s_58;
    _zz_io_s_61 <= _zz_io_s_60[56:0];
    _zz_io_s_62 <= _zz_io_s_60[57];
  end


endmodule

module FineReduction (
  input      [377:0]  io_a,
  output     [376:0]  io_r,
  input               clk,
  input               resetn
);

  wire       [378:0]  singleAdd_add_io_s;
  wire       [376:0]  _zz__zz_io_r;
  wire       [376:0]  _zz__zz_io_r_1;
  reg        [377:0]  io_a_delay_1;
  reg        [377:0]  io_a_delay_2;
  reg        [377:0]  io_a_delay_3;
  reg        [377:0]  io_a_delay_4;
  reg        [377:0]  io_a_delay_5;
  reg        [377:0]  singleAdd_a;
  reg        [376:0]  _zz_io_r;

  assign _zz__zz_io_r = singleAdd_a[376:0];
  assign _zz__zz_io_r_1 = singleAdd_add_io_s[376:0];
  BADD_1 singleAdd_add (
    .io_a   (io_a[377:0]                                                                                         ), //i
    .io_b   (378'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001), //i
    .io_c   (1'b1                                                                                                ), //i
    .io_s   (singleAdd_add_io_s[378:0]                                                                           ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  assign io_r = _zz_io_r;
  always @(posedge clk) begin
    io_a_delay_1 <= io_a;
    io_a_delay_2 <= io_a_delay_1;
    io_a_delay_3 <= io_a_delay_2;
    io_a_delay_4 <= io_a_delay_3;
    io_a_delay_5 <= io_a_delay_4;
    singleAdd_a <= io_a_delay_5;
    _zz_io_r <= (singleAdd_add_io_s[377] ? _zz__zz_io_r : _zz__zz_io_r_1);
  end


endmodule

//MADD_7 replaced by MADD_4

//MADD_6 replaced by MADD_4

//MADD_5 replaced by MADD_4

module MADD_4 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  output     [376:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [377:0]  add_io_s;
  wire       [376:0]  reduction_io_r;

  BADD_5 add (
    .io_a   (io_a[376:0]    ), //i
    .io_b   (io_b[376:0]    ), //i
    .io_c   (1'b1           ), //i
    .io_s   (add_io_s[377:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  FineReduction_26 reduction (
    .io_a   (add_io_s[377:0]      ), //i
    .io_r   (reduction_io_r[376:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign io_s = reduction_io_r;

endmodule

//MADD_3 replaced by MADD

//MADD_2 replaced by MADD

//MADD_1 replaced by MADD

module MADD (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  output     [376:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [377:0]  add_io_s;
  wire       [376:0]  reduction_io_r;

  BADD_9 add (
    .io_a   (io_a[376:0]    ), //i
    .io_b   (io_b[376:0]    ), //i
    .io_c   (1'b0           ), //i
    .io_s   (add_io_s[377:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  FineReduction_8 reduction (
    .io_a   (add_io_s[377:0]      ), //i
    .io_r   (reduction_io_r[376:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign io_s = reduction_io_r;

endmodule

//KaratsubaMMUL_8 replaced by KaratsubaMMUL

//KaratsubaMMUL_7 replaced by KaratsubaMMUL

//KaratsubaMMUL_6 replaced by KaratsubaMMUL

//KaratsubaMMUL_5 replaced by KaratsubaMMUL

//KaratsubaMMUL_4 replaced by KaratsubaMMUL

//KaratsubaMMUL_3 replaced by KaratsubaMMUL

//KaratsubaMMUL_2 replaced by KaratsubaMMUL

//KaratsubaMMUL_1 replaced by KaratsubaMMUL

module KaratsubaMMUL (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  output     [376:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [377:0]  useBarrett_cMul1_io_a;
  wire       [377:0]  useBarrett_cMul2_io_a;
  wire       [378:0]  useBarrett_reduction_io_a;
  wire       [753:0]  useBarrett_mul_io_p;
  wire       [755:0]  useBarrett_cMul1_io_p;
  wire       [378:0]  useBarrett_cMul2_io_p;
  wire       [379:0]  useBarrett_sub_io_s;
  wire       [376:0]  useBarrett_reduction_io_r;
  reg        [378:0]  _zz_io_a;
  reg        [378:0]  _zz_io_a_1;
  reg        [378:0]  _zz_io_a_2;
  reg        [378:0]  _zz_io_a_3;
  reg        [378:0]  _zz_io_a_4;
  reg        [378:0]  _zz_io_a_5;
  reg        [378:0]  _zz_io_a_6;
  reg        [378:0]  _zz_io_a_7;
  reg        [378:0]  _zz_io_a_8;
  reg        [378:0]  _zz_io_a_9;
  reg        [378:0]  _zz_io_a_10;
  reg        [378:0]  _zz_io_a_11;
  reg        [378:0]  _zz_io_a_12;
  reg        [378:0]  _zz_io_a_13;
  reg        [378:0]  _zz_io_a_14;
  reg        [378:0]  _zz_io_a_15;
  reg        [378:0]  _zz_io_a_16;
  reg        [378:0]  _zz_io_a_17;
  reg        [378:0]  _zz_io_a_18;
  reg        [378:0]  _zz_io_a_19;
  reg        [378:0]  _zz_io_a_20;
  reg        [378:0]  _zz_io_a_21;
  reg        [378:0]  _zz_io_a_22;
  reg        [378:0]  _zz_io_a_23;
  reg        [378:0]  _zz_io_a_24;
  reg        [378:0]  _zz_io_a_25;
  reg        [378:0]  _zz_io_a_26;
  reg        [378:0]  _zz_io_a_27;
  reg        [378:0]  _zz_io_a_28;
  reg        [378:0]  _zz_io_a_29;
  reg        [378:0]  _zz_io_a_30;
  reg        [378:0]  _zz_io_a_31;
  reg        [378:0]  _zz_io_a_32;
  reg        [378:0]  _zz_io_a_33;
  reg        [378:0]  _zz_io_a_34;
  reg        [378:0]  _zz_io_a_35;
  reg        [378:0]  _zz_io_a_36;
  reg        [378:0]  _zz_io_a_37;
  reg        [378:0]  _zz_io_a_38;
  reg        [378:0]  _zz_io_a_39;
  reg        [378:0]  _zz_io_a_40;

  KaratsubaMUL_16 useBarrett_mul (
    .io_a   (io_a[376:0]               ), //i
    .io_b   (io_b[376:0]               ), //i
    .io_p   (useBarrett_mul_io_p[753:0]), //o
    .clk    (clk                       ), //i
    .resetn (resetn                    )  //i
  );
  KaratsubaMUL_17 useBarrett_cMul1 (
    .io_a   (useBarrett_cMul1_io_a[377:0]                                                                        ), //i
    .io_b   (378'h261508d0cc4060e976c3ca0582ef4f73bbad0de6776b1a06af2d488d85a6d02d0ed687789c42a591f9fd58c5e4daffc), //i
    .io_p   (useBarrett_cMul1_io_p[755:0]                                                                        ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  BCMUL_8 useBarrett_cMul2 (
    .io_a   (useBarrett_cMul2_io_a[377:0]), //i
    .io_p   (useBarrett_cMul2_io_p[378:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_18 useBarrett_sub (
    .io_a   (_zz_io_a_40[378:0]          ), //i
    .io_b   (useBarrett_cMul2_io_p[378:0]), //i
    .io_c   (1'b1                        ), //i
    .io_s   (useBarrett_sub_io_s[379:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  FineReduction_17 useBarrett_reduction (
    .io_a   (useBarrett_reduction_io_a[378:0]), //i
    .io_r   (useBarrett_reduction_io_r[376:0]), //o
    .clk    (clk                             ), //i
    .resetn (resetn                          )  //i
  );
  assign useBarrett_cMul1_io_a = useBarrett_mul_io_p[753 : 376];
  assign useBarrett_cMul2_io_a = useBarrett_cMul1_io_p[755 : 378];
  assign useBarrett_reduction_io_a = useBarrett_sub_io_s[378:0];
  assign io_p = useBarrett_reduction_io_r;
  always @(posedge clk) begin
    _zz_io_a <= useBarrett_mul_io_p[378:0];
    _zz_io_a_1 <= _zz_io_a;
    _zz_io_a_2 <= _zz_io_a_1;
    _zz_io_a_3 <= _zz_io_a_2;
    _zz_io_a_4 <= _zz_io_a_3;
    _zz_io_a_5 <= _zz_io_a_4;
    _zz_io_a_6 <= _zz_io_a_5;
    _zz_io_a_7 <= _zz_io_a_6;
    _zz_io_a_8 <= _zz_io_a_7;
    _zz_io_a_9 <= _zz_io_a_8;
    _zz_io_a_10 <= _zz_io_a_9;
    _zz_io_a_11 <= _zz_io_a_10;
    _zz_io_a_12 <= _zz_io_a_11;
    _zz_io_a_13 <= _zz_io_a_12;
    _zz_io_a_14 <= _zz_io_a_13;
    _zz_io_a_15 <= _zz_io_a_14;
    _zz_io_a_16 <= _zz_io_a_15;
    _zz_io_a_17 <= _zz_io_a_16;
    _zz_io_a_18 <= _zz_io_a_17;
    _zz_io_a_19 <= _zz_io_a_18;
    _zz_io_a_20 <= _zz_io_a_19;
    _zz_io_a_21 <= _zz_io_a_20;
    _zz_io_a_22 <= _zz_io_a_21;
    _zz_io_a_23 <= _zz_io_a_22;
    _zz_io_a_24 <= _zz_io_a_23;
    _zz_io_a_25 <= _zz_io_a_24;
    _zz_io_a_26 <= _zz_io_a_25;
    _zz_io_a_27 <= _zz_io_a_26;
    _zz_io_a_28 <= _zz_io_a_27;
    _zz_io_a_29 <= _zz_io_a_28;
    _zz_io_a_30 <= _zz_io_a_29;
    _zz_io_a_31 <= _zz_io_a_30;
    _zz_io_a_32 <= _zz_io_a_31;
    _zz_io_a_33 <= _zz_io_a_32;
    _zz_io_a_34 <= _zz_io_a_33;
    _zz_io_a_35 <= _zz_io_a_34;
    _zz_io_a_36 <= _zz_io_a_35;
    _zz_io_a_37 <= _zz_io_a_36;
    _zz_io_a_38 <= _zz_io_a_37;
    _zz_io_a_39 <= _zz_io_a_38;
    _zz_io_a_40 <= _zz_io_a_39;
  end


endmodule

module SDPRAM (
  input               io_we,
  input      [7:0]    io_wAddress,
  input      [376:0]  io_wData_a_X,
  input      [376:0]  io_wData_a_Y,
  input      [376:0]  io_wData_a_Z,
  input      [376:0]  io_wData_a_T,
  input      [376:0]  io_wData_b_X,
  input      [376:0]  io_wData_b_Y,
  input      [376:0]  io_wData_b_Z,
  input      [376:0]  io_wData_b_T,
  input      [16:0]   io_wData_address,
  input               io_re,
  input      [7:0]    io_rAddress,
  output     [376:0]  io_rData_a_X,
  output     [376:0]  io_rData_a_Y,
  output     [376:0]  io_rData_a_Z,
  output     [376:0]  io_rData_a_T,
  output     [376:0]  io_rData_b_X,
  output     [376:0]  io_rData_b_Y,
  output     [376:0]  io_rData_b_Z,
  output     [376:0]  io_rData_b_T,
  output     [16:0]   io_rData_address,
  input               clk,
  input               resetn
);

  wire       [3032:0] ram_doutb;
  reg        [7:0]    io_wAddress_regNext;
  reg        [3032:0] _zz_dina;
  reg                 io_we_regNext;
  reg        [7:0]    io_rAddress_regNext;
  reg                 io_re_regNext;
  wire       [1507:0] _zz_io_rData_a_X;
  wire       [1507:0] _zz_io_rData_b_X;

  xpm_memory_sdpram #(
    .ADDR_WIDTH_A(8),
    .ADDR_WIDTH_B(8),
    .AUTO_SLEEP_TIME(0),
    .BYTE_WRITE_WIDTH_A(3033),
    .CASCADE_HEIGHT(0),
    .CLOCKING_MODE("common_clock"),
    .ECC_MODE("no_ecc"),
    .MEMORY_INIT_FILE("none"),
    .MEMORY_INIT_PARAM("0"),
    .MEMORY_OPTIMIZATION("true"),
    .MEMORY_PRIMITIVE("auto"),
    .MEMORY_SIZE(776448),
    .MESSAGE_CONTROL(0),
    .READ_DATA_WIDTH_B(3033),
    .READ_LATENCY_B(3),
    .READ_RESET_VALUE_B("0"),
    .RST_MODE_A("SYNC"),
    .RST_MODE_B("SYNC"),
    .SIM_ASSERT_CHK(0),
    .USE_EMBEDDED_CONSTRAINT(0),
    .USE_MEM_INIT(1),
    .WAKEUP_TIME("disable_sleep"),
    .WRITE_DATA_WIDTH_A(3033),
    .WRITE_MODE_B("read_first"),
    .WRITE_PROTECT(1)
  ) ram (
    .addra          (io_wAddress_regNext[7:0]), //i
    .addrb          (io_rAddress_regNext[7:0]), //i
    .dina           (_zz_dina[3032:0]        ), //i
    .doutb          (ram_doutb[3032:0]       ), //o
    .enb            (io_re_regNext           ), //i
    .wea            (io_we_regNext           ), //i
    .clka           (clk                     ), //i
    .clkb           (clk                     ), //i
    .ena            (1'b1                    ), //i
    .injectdbiterra (1'b0                    ), //i
    .injectsbiterra (1'b0                    ), //i
    .regceb         (1'b1                    ), //i
    .rstb           (1'b0                    ), //i
    .sleep          (1'b0                    )  //i
  );
  assign _zz_io_rData_a_X = ram_doutb[1507 : 0];
  assign io_rData_a_X = _zz_io_rData_a_X[376 : 0];
  assign io_rData_a_Y = _zz_io_rData_a_X[753 : 377];
  assign io_rData_a_Z = _zz_io_rData_a_X[1130 : 754];
  assign io_rData_a_T = _zz_io_rData_a_X[1507 : 1131];
  assign _zz_io_rData_b_X = ram_doutb[3015 : 1508];
  assign io_rData_b_X = _zz_io_rData_b_X[376 : 0];
  assign io_rData_b_Y = _zz_io_rData_b_X[753 : 377];
  assign io_rData_b_Z = _zz_io_rData_b_X[1130 : 754];
  assign io_rData_b_T = _zz_io_rData_b_X[1507 : 1131];
  assign io_rData_address = ram_doutb[3032 : 3016];
  always @(posedge clk) begin
    io_wAddress_regNext <= io_wAddress;
    _zz_dina <= {io_wData_address,{{io_wData_b_T,{io_wData_b_Z,{io_wData_b_Y,io_wData_b_X}}},{io_wData_a_T,{io_wData_a_Z,{io_wData_a_Y,io_wData_a_X}}}}};
    io_we_regNext <= io_we;
    io_rAddress_regNext <= io_rAddress;
    io_re_regNext <= io_re;
  end


endmodule

module TDPRAM (
  input               io_we_0,
  input               io_we_1,
  input      [16:0]   io_address_0,
  input      [16:0]   io_address_1,
  input      [376:0]  io_wData_0_X,
  input      [376:0]  io_wData_0_Y,
  input      [376:0]  io_wData_0_Z,
  input      [376:0]  io_wData_0_T,
  input      [376:0]  io_wData_1_X,
  input      [376:0]  io_wData_1_Y,
  input      [376:0]  io_wData_1_Z,
  input      [376:0]  io_wData_1_T,
  input               io_ce_0,
  input               io_ce_1,
  output     [376:0]  io_rData_0_X,
  output     [376:0]  io_rData_0_Y,
  output     [376:0]  io_rData_0_Z,
  output     [376:0]  io_rData_0_T,
  output     [376:0]  io_rData_1_X,
  output     [376:0]  io_rData_1_Y,
  output     [376:0]  io_rData_1_Z,
  output     [376:0]  io_rData_1_T,
  input               clk,
  input               resetn
);

  wire       [1507:0] ram_douta;
  wire       [1507:0] ram_doutb;
  reg        [16:0]   io_address_0_regNext;
  reg        [1507:0] _zz_dina;
  reg                 io_ce_0_regNext;
  reg                 io_we_0_regNext;
  reg        [16:0]   io_address_1_regNext;
  reg        [1507:0] _zz_dinb;
  reg                 io_ce_1_regNext;
  reg                 io_we_1_regNext;

  xpm_memory_tdpram #(
    .ADDR_WIDTH_A(17),
    .ADDR_WIDTH_B(17),
    .AUTO_SLEEP_TIME(0),
    .BYTE_WRITE_WIDTH_A(1508),
    .BYTE_WRITE_WIDTH_B(1508),
    .CASCADE_HEIGHT(0),
    .CLOCKING_MODE("common_clock"),
    .ECC_MODE("no_ecc"),
    .MEMORY_INIT_FILE("none"),
    .MEMORY_INIT_PARAM("0"),
    .MEMORY_OPTIMIZATION("true"),
    .MEMORY_PRIMITIVE("ultra"),
    .MEMORY_SIZE(123535360),
    .MESSAGE_CONTROL(0),
    .READ_DATA_WIDTH_A(1508),
    .READ_DATA_WIDTH_B(1508),
    .READ_LATENCY_A(28),
    .READ_LATENCY_B(28),
    .READ_RESET_VALUE_A("0"),
    .READ_RESET_VALUE_B("0"),
    .RST_MODE_A("SYNC"),
    .RST_MODE_B("SYNC"),
    .SIM_ASSERT_CHK(0),
    .USE_EMBEDDED_CONSTRAINT(0),
    .USE_MEM_INIT(1),
    .USE_MEM_INIT_MMI(0),
    .WAKEUP_TIME("disable_sleep"),
    .WRITE_DATA_WIDTH_A(1508),
    .WRITE_DATA_WIDTH_B(1508),
    .WRITE_MODE_A("no_change"),
    .WRITE_MODE_B("no_change"),
    .WRITE_PROTECT(1)
  ) ram (
    .addra          (io_address_0_regNext[16:0]), //i
    .addrb          (io_address_1_regNext[16:0]), //i
    .dina           (_zz_dina[1507:0]          ), //i
    .dinb           (_zz_dinb[1507:0]          ), //i
    .douta          (ram_douta[1507:0]         ), //o
    .doutb          (ram_doutb[1507:0]         ), //o
    .ena            (io_ce_0_regNext           ), //i
    .enb            (io_ce_1_regNext           ), //i
    .wea            (io_we_0_regNext           ), //i
    .web            (io_we_1_regNext           ), //i
    .clka           (clk                       ), //i
    .clkb           (clk                       ), //i
    .injectdbiterra (1'b0                      ), //i
    .injectdbiterrb (1'b0                      ), //i
    .injectsbiterra (1'b0                      ), //i
    .injectsbiterrb (1'b0                      ), //i
    .regcea         (1'b1                      ), //i
    .regceb         (1'b1                      ), //i
    .rsta           (1'b0                      ), //i
    .rstb           (1'b0                      ), //i
    .sleep          (1'b0                      )  //i
  );
  assign io_rData_0_X = ram_douta[376 : 0];
  assign io_rData_0_Y = ram_douta[753 : 377];
  assign io_rData_0_Z = ram_douta[1130 : 754];
  assign io_rData_0_T = ram_douta[1507 : 1131];
  assign io_rData_1_X = ram_doutb[376 : 0];
  assign io_rData_1_Y = ram_doutb[753 : 377];
  assign io_rData_1_Z = ram_doutb[1130 : 754];
  assign io_rData_1_T = ram_doutb[1507 : 1131];
  always @(posedge clk) begin
    io_address_0_regNext <= io_address_0;
    _zz_dina <= {io_wData_0_T,{io_wData_0_Z,{io_wData_0_Y,io_wData_0_X}}};
    io_ce_0_regNext <= io_ce_0;
    io_we_0_regNext <= io_we_0;
    io_address_1_regNext <= io_address_1;
    _zz_dinb <= {io_wData_1_T,{io_wData_1_Z,{io_wData_1_Y,io_wData_1_X}}};
    io_ce_1_regNext <= io_ce_1;
    io_we_1_regNext <= io_we_1;
  end


endmodule

//SDPRAM_4 replaced by SDPRAM_1

//SDPRAM_3 replaced by SDPRAM_1

//SDPRAM_2 replaced by SDPRAM_1

module SDPRAM_1 (
  input               io_we,
  input      [16:0]   io_wAddress,
  input               io_wData,
  input               io_re,
  input      [16:0]   io_rAddress,
  output              io_rData,
  input               clk,
  input               resetn
);

  wire       [0:0]    ram_doutb;
  reg        [16:0]   io_wAddress_regNext;
  reg        [0:0]    _zz_dina;
  reg                 io_we_regNext;
  reg        [16:0]   io_rAddress_regNext;
  reg                 io_re_regNext;

  xpm_memory_sdpram #(
    .ADDR_WIDTH_A(17),
    .ADDR_WIDTH_B(17),
    .AUTO_SLEEP_TIME(0),
    .BYTE_WRITE_WIDTH_A(1),
    .CASCADE_HEIGHT(0),
    .CLOCKING_MODE("common_clock"),
    .ECC_MODE("no_ecc"),
    .MEMORY_INIT_FILE("none"),
    .MEMORY_INIT_PARAM("0"),
    .MEMORY_OPTIMIZATION("true"),
    .MEMORY_PRIMITIVE("auto"),
    .MEMORY_SIZE(81920),
    .MESSAGE_CONTROL(0),
    .READ_DATA_WIDTH_B(1),
    .READ_LATENCY_B(2),
    .READ_RESET_VALUE_B("0"),
    .RST_MODE_A("SYNC"),
    .RST_MODE_B("SYNC"),
    .SIM_ASSERT_CHK(0),
    .USE_EMBEDDED_CONSTRAINT(0),
    .USE_MEM_INIT(1),
    .WAKEUP_TIME("disable_sleep"),
    .WRITE_DATA_WIDTH_A(1),
    .WRITE_MODE_B("read_first"),
    .WRITE_PROTECT(1)
  ) ram (
    .addra          (io_wAddress_regNext[16:0]), //i
    .addrb          (io_rAddress_regNext[16:0]), //i
    .dina           (_zz_dina                 ), //i
    .doutb          (ram_doutb                ), //o
    .enb            (io_re_regNext            ), //i
    .wea            (io_we_regNext            ), //i
    .clka           (clk                      ), //i
    .clkb           (clk                      ), //i
    .ena            (1'b1                     ), //i
    .injectdbiterra (1'b0                     ), //i
    .injectsbiterra (1'b0                     ), //i
    .regceb         (1'b1                     ), //i
    .rstb           (1'b0                     ), //i
    .sleep          (1'b0                     )  //i
  );
  assign io_rData = ram_doutb[0];
  always @(posedge clk) begin
    io_wAddress_regNext <= io_wAddress;
    _zz_dina <= io_wData;
    io_we_regNext <= io_we;
    io_rAddress_regNext <= io_rAddress;
    io_re_regNext <= io_re;
  end


endmodule

module BADD_1 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  input               io_c,
  output reg [378:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [377:0]  _zz__zz_io_s_1;
  wire       [64:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [377:0]  _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_10;
  wire       [64:0]   _zz__zz_io_s_10_1;
  wire       [0:0]    _zz__zz_io_s_10_2;
  wire       [377:0]  _zz__zz_io_s_19;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [377:0]  _zz__zz_io_s_30;
  wire       [64:0]   _zz__zz_io_s_33;
  wire       [64:0]   _zz__zz_io_s_33_1;
  wire       [0:0]    _zz__zz_io_s_33_2;
  wire       [377:0]  _zz__zz_io_s_42;
  wire       [64:0]   _zz__zz_io_s_46;
  wire       [64:0]   _zz__zz_io_s_46_1;
  wire       [0:0]    _zz__zz_io_s_46_2;
  wire       [377:0]  _zz__zz_io_s_55;
  wire       [58:0]   _zz__zz_io_s_60;
  wire       [58:0]   _zz__zz_io_s_60_1;
  wire       [0:0]    _zz__zz_io_s_60_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  wire       [64:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg                 _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg        [63:0]   _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg        [63:0]   _zz_io_s_25;
  reg                 _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg        [63:0]   _zz_io_s_29;
  reg        [63:0]   _zz_io_s_30;
  reg        [63:0]   _zz_io_s_31;
  reg        [63:0]   _zz_io_s_32;
  wire       [64:0]   _zz_io_s_33;
  reg        [63:0]   _zz_io_s_34;
  reg        [63:0]   _zz_io_s_35;
  reg        [63:0]   _zz_io_s_36;
  reg                 _zz_io_s_37;
  reg        [63:0]   _zz_io_s_38;
  reg        [63:0]   _zz_io_s_39;
  reg        [63:0]   _zz_io_s_40;
  reg        [63:0]   _zz_io_s_41;
  reg        [63:0]   _zz_io_s_42;
  reg        [63:0]   _zz_io_s_43;
  reg        [63:0]   _zz_io_s_44;
  reg        [63:0]   _zz_io_s_45;
  wire       [64:0]   _zz_io_s_46;
  reg        [63:0]   _zz_io_s_47;
  reg        [63:0]   _zz_io_s_48;
  reg                 _zz_io_s_49;
  reg        [57:0]   _zz_io_s_50;
  reg        [57:0]   _zz_io_s_51;
  reg        [57:0]   _zz_io_s_52;
  reg        [57:0]   _zz_io_s_53;
  reg        [57:0]   _zz_io_s_54;
  reg        [57:0]   _zz_io_s_55;
  reg        [57:0]   _zz_io_s_56;
  reg        [57:0]   _zz_io_s_57;
  reg        [57:0]   _zz_io_s_58;
  reg        [57:0]   _zz_io_s_59;
  wire       [58:0]   _zz_io_s_60;
  reg        [57:0]   _zz_io_s_61;
  reg                 _zz_io_s_62;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,_zz__zz_io_s_1[63 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {64'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_9 = (~ io_b);
  assign _zz__zz_io_s_10 = ({1'b0,_zz_io_s_8} + {1'b0,_zz_io_s_9});
  assign _zz__zz_io_s_10_2 = _zz_io_s_7;
  assign _zz__zz_io_s_10_1 = {64'd0, _zz__zz_io_s_10_2};
  assign _zz__zz_io_s_19 = (~ io_b);
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_18} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_16;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_30 = (~ io_b);
  assign _zz__zz_io_s_33 = ({1'b0,_zz_io_s_29} + {1'b0,_zz_io_s_32});
  assign _zz__zz_io_s_33_2 = _zz_io_s_26;
  assign _zz__zz_io_s_33_1 = {64'd0, _zz__zz_io_s_33_2};
  assign _zz__zz_io_s_42 = (~ io_b);
  assign _zz__zz_io_s_46 = ({1'b0,_zz_io_s_41} + {1'b0,_zz_io_s_45});
  assign _zz__zz_io_s_46_2 = _zz_io_s_37;
  assign _zz__zz_io_s_46_1 = {64'd0, _zz__zz_io_s_46_2};
  assign _zz__zz_io_s_55 = (~ io_b);
  assign _zz__zz_io_s_60 = ({1'b0,_zz_io_s_54} + {1'b0,_zz_io_s_59});
  assign _zz__zz_io_s_60_2 = _zz_io_s_49;
  assign _zz__zz_io_s_60_1 = {58'd0, _zz__zz_io_s_60_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_6;
    io_s[127 : 64] = _zz_io_s_15;
    io_s[191 : 128] = _zz_io_s_25;
    io_s[255 : 192] = _zz_io_s_36;
    io_s[319 : 256] = _zz_io_s_48;
    io_s[377 : 320] = _zz_io_s_61;
    io_s[378] = (! _zz_io_s_62);
  end

  assign _zz_io_s_10 = (_zz__zz_io_s_10 + _zz__zz_io_s_10_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_33 = (_zz__zz_io_s_33 + _zz__zz_io_s_33_1);
  assign _zz_io_s_46 = (_zz__zz_io_s_46 + _zz__zz_io_s_46_1);
  assign _zz_io_s_60 = (_zz__zz_io_s_60 + _zz__zz_io_s_60_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= _zz_io_s[64];
    _zz_io_s_8 <= io_a[127 : 64];
    _zz_io_s_9 <= _zz__zz_io_s_9[127 : 64];
    _zz_io_s_11 <= _zz_io_s_10[63:0];
    _zz_io_s_12 <= _zz_io_s_11;
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= _zz_io_s_10[64];
    _zz_io_s_17 <= io_a[191 : 128];
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= _zz__zz_io_s_19[191 : 128];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_22;
    _zz_io_s_24 <= _zz_io_s_23;
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_21[64];
    _zz_io_s_27 <= io_a[255 : 192];
    _zz_io_s_28 <= _zz_io_s_27;
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz__zz_io_s_30[255 : 192];
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_32 <= _zz_io_s_31;
    _zz_io_s_34 <= _zz_io_s_33[63:0];
    _zz_io_s_35 <= _zz_io_s_34;
    _zz_io_s_36 <= _zz_io_s_35;
    _zz_io_s_37 <= _zz_io_s_33[64];
    _zz_io_s_38 <= io_a[319 : 256];
    _zz_io_s_39 <= _zz_io_s_38;
    _zz_io_s_40 <= _zz_io_s_39;
    _zz_io_s_41 <= _zz_io_s_40;
    _zz_io_s_42 <= _zz__zz_io_s_42[319 : 256];
    _zz_io_s_43 <= _zz_io_s_42;
    _zz_io_s_44 <= _zz_io_s_43;
    _zz_io_s_45 <= _zz_io_s_44;
    _zz_io_s_47 <= _zz_io_s_46[63:0];
    _zz_io_s_48 <= _zz_io_s_47;
    _zz_io_s_49 <= _zz_io_s_46[64];
    _zz_io_s_50 <= io_a[377 : 320];
    _zz_io_s_51 <= _zz_io_s_50;
    _zz_io_s_52 <= _zz_io_s_51;
    _zz_io_s_53 <= _zz_io_s_52;
    _zz_io_s_54 <= _zz_io_s_53;
    _zz_io_s_55 <= _zz__zz_io_s_55[377 : 320];
    _zz_io_s_56 <= _zz_io_s_55;
    _zz_io_s_57 <= _zz_io_s_56;
    _zz_io_s_58 <= _zz_io_s_57;
    _zz_io_s_59 <= _zz_io_s_58;
    _zz_io_s_61 <= _zz_io_s_60[57:0];
    _zz_io_s_62 <= _zz_io_s_60[58];
  end


endmodule

//FineReduction_1 replaced by FineReduction_26

//BADD_2 replaced by BADD_5

//FineReduction_2 replaced by FineReduction_26

//BADD_3 replaced by BADD_5

//FineReduction_3 replaced by FineReduction_26

//BADD_4 replaced by BADD_5

//FineReduction_4 replaced by FineReduction_26

module BADD_5 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  input               io_c,
  output reg [377:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [376:0]  _zz__zz_io_s_1;
  wire       [64:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [376:0]  _zz__zz_io_s_4;
  wire       [64:0]   _zz__zz_io_s_5;
  wire       [64:0]   _zz__zz_io_s_5_1;
  wire       [0:0]    _zz__zz_io_s_5_2;
  wire       [376:0]  _zz__zz_io_s_10;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [376:0]  _zz__zz_io_s_18;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [376:0]  _zz__zz_io_s_28;
  wire       [64:0]   _zz__zz_io_s_32;
  wire       [64:0]   _zz__zz_io_s_32_1;
  wire       [0:0]    _zz__zz_io_s_32_2;
  wire       [376:0]  _zz__zz_io_s_40;
  wire       [57:0]   _zz__zz_io_s_45;
  wire       [57:0]   _zz__zz_io_s_45_1;
  wire       [0:0]    _zz__zz_io_s_45_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  wire       [64:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg        [63:0]   _zz_io_s_25;
  reg        [63:0]   _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg        [63:0]   _zz_io_s_29;
  reg        [63:0]   _zz_io_s_30;
  reg        [63:0]   _zz_io_s_31;
  wire       [64:0]   _zz_io_s_32;
  reg        [63:0]   _zz_io_s_33;
  reg                 _zz_io_s_34;
  reg        [56:0]   _zz_io_s_35;
  reg        [56:0]   _zz_io_s_36;
  reg        [56:0]   _zz_io_s_37;
  reg        [56:0]   _zz_io_s_38;
  reg        [56:0]   _zz_io_s_39;
  reg        [56:0]   _zz_io_s_40;
  reg        [56:0]   _zz_io_s_41;
  reg        [56:0]   _zz_io_s_42;
  reg        [56:0]   _zz_io_s_43;
  reg        [56:0]   _zz_io_s_44;
  wire       [57:0]   _zz_io_s_45;
  reg        [56:0]   _zz_io_s_46;
  reg                 _zz_io_s_47;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,_zz__zz_io_s_1[63 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {64'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_4 = (~ io_b);
  assign _zz__zz_io_s_5 = ({1'b0,_zz_io_s_3} + {1'b0,_zz_io_s_4});
  assign _zz__zz_io_s_5_2 = _zz_io_s_2;
  assign _zz__zz_io_s_5_1 = {64'd0, _zz__zz_io_s_5_2};
  assign _zz__zz_io_s_10 = (~ io_b);
  assign _zz__zz_io_s_12 = ({1'b0,_zz_io_s_9} + {1'b0,_zz_io_s_11});
  assign _zz__zz_io_s_12_2 = _zz_io_s_7;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_18 = (~ io_b);
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_17} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_14;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_28 = (~ io_b);
  assign _zz__zz_io_s_32 = ({1'b0,_zz_io_s_27} + {1'b0,_zz_io_s_31});
  assign _zz__zz_io_s_32_2 = _zz_io_s_23;
  assign _zz__zz_io_s_32_1 = {64'd0, _zz__zz_io_s_32_2};
  assign _zz__zz_io_s_40 = (~ io_b);
  assign _zz__zz_io_s_45 = ({1'b0,_zz_io_s_39} + {1'b0,_zz_io_s_44});
  assign _zz__zz_io_s_45_2 = _zz_io_s_34;
  assign _zz__zz_io_s_45_1 = {57'd0, _zz__zz_io_s_45_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_1;
    io_s[127 : 64] = _zz_io_s_6;
    io_s[191 : 128] = _zz_io_s_13;
    io_s[255 : 192] = _zz_io_s_22;
    io_s[319 : 256] = _zz_io_s_33;
    io_s[376 : 320] = _zz_io_s_46;
    io_s[377] = (! _zz_io_s_47);
  end

  assign _zz_io_s_5 = (_zz__zz_io_s_5 + _zz__zz_io_s_5_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_32 = (_zz__zz_io_s_32 + _zz__zz_io_s_32_1);
  assign _zz_io_s_45 = (_zz__zz_io_s_45 + _zz__zz_io_s_45_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s[64];
    _zz_io_s_3 <= io_a[127 : 64];
    _zz_io_s_4 <= _zz__zz_io_s_4[127 : 64];
    _zz_io_s_6 <= _zz_io_s_5[63:0];
    _zz_io_s_7 <= _zz_io_s_5[64];
    _zz_io_s_8 <= io_a[191 : 128];
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz__zz_io_s_10[191 : 128];
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_15 <= io_a[255 : 192];
    _zz_io_s_16 <= _zz_io_s_15;
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz__zz_io_s_18[255 : 192];
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_21[64];
    _zz_io_s_24 <= io_a[319 : 256];
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_25;
    _zz_io_s_27 <= _zz_io_s_26;
    _zz_io_s_28 <= _zz__zz_io_s_28[319 : 256];
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz_io_s_29;
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_33 <= _zz_io_s_32[63:0];
    _zz_io_s_34 <= _zz_io_s_32[64];
    _zz_io_s_35 <= io_a[376 : 320];
    _zz_io_s_36 <= _zz_io_s_35;
    _zz_io_s_37 <= _zz_io_s_36;
    _zz_io_s_38 <= _zz_io_s_37;
    _zz_io_s_39 <= _zz_io_s_38;
    _zz_io_s_40 <= _zz__zz_io_s_40[376 : 320];
    _zz_io_s_41 <= _zz_io_s_40;
    _zz_io_s_42 <= _zz_io_s_41;
    _zz_io_s_43 <= _zz_io_s_42;
    _zz_io_s_44 <= _zz_io_s_43;
    _zz_io_s_46 <= _zz_io_s_45[56:0];
    _zz_io_s_47 <= _zz_io_s_45[57];
  end


endmodule

//FineReduction_5 replaced by FineReduction_8

//BADD_6 replaced by BADD_9

//FineReduction_6 replaced by FineReduction_8

//BADD_7 replaced by BADD_9

//FineReduction_7 replaced by FineReduction_8

//BADD_8 replaced by BADD_9

module FineReduction_8 (
  input      [377:0]  io_a,
  output     [376:0]  io_r,
  input               clk,
  input               resetn
);

  wire       [378:0]  singleAdd_add_io_s;
  wire       [376:0]  _zz__zz_io_r;
  wire       [376:0]  _zz__zz_io_r_1;
  reg        [63:0]   _zz_singleAdd_a;
  reg        [63:0]   _zz_singleAdd_a_1;
  reg        [63:0]   _zz_singleAdd_a_2;
  reg        [63:0]   _zz_singleAdd_a_3;
  reg        [63:0]   _zz_singleAdd_a_4;
  reg        [63:0]   _zz_singleAdd_a_5;
  reg        [63:0]   _zz_singleAdd_a_6;
  reg        [63:0]   _zz_singleAdd_a_7;
  reg        [63:0]   _zz_singleAdd_a_8;
  reg        [63:0]   _zz_singleAdd_a_9;
  reg        [63:0]   _zz_singleAdd_a_10;
  reg        [63:0]   _zz_singleAdd_a_11;
  reg        [63:0]   _zz_singleAdd_a_12;
  reg        [63:0]   _zz_singleAdd_a_13;
  reg        [63:0]   _zz_singleAdd_a_14;
  reg        [63:0]   _zz_singleAdd_a_15;
  reg        [63:0]   _zz_singleAdd_a_16;
  reg        [63:0]   _zz_singleAdd_a_17;
  reg        [63:0]   _zz_singleAdd_a_18;
  reg        [63:0]   _zz_singleAdd_a_19;
  reg        [57:0]   _zz_singleAdd_a_20;
  wire       [377:0]  singleAdd_a;
  reg        [376:0]  _zz_io_r;

  assign _zz__zz_io_r = singleAdd_a[376:0];
  assign _zz__zz_io_r_1 = singleAdd_add_io_s[376:0];
  BADD_26 singleAdd_add (
    .io_a   (io_a[377:0]                                                                                         ), //i
    .io_b   (378'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001), //i
    .io_c   (1'b1                                                                                                ), //i
    .io_s   (singleAdd_add_io_s[378:0]                                                                           ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  assign singleAdd_a = {_zz_singleAdd_a_20,{_zz_singleAdd_a_19,{_zz_singleAdd_a_17,{_zz_singleAdd_a_14,{_zz_singleAdd_a_10,_zz_singleAdd_a_5}}}}};
  assign io_r = _zz_io_r;
  always @(posedge clk) begin
    _zz_singleAdd_a <= io_a[63 : 0];
    _zz_singleAdd_a_1 <= _zz_singleAdd_a;
    _zz_singleAdd_a_2 <= _zz_singleAdd_a_1;
    _zz_singleAdd_a_3 <= _zz_singleAdd_a_2;
    _zz_singleAdd_a_4 <= _zz_singleAdd_a_3;
    _zz_singleAdd_a_5 <= _zz_singleAdd_a_4;
    _zz_singleAdd_a_6 <= io_a[127 : 64];
    _zz_singleAdd_a_7 <= _zz_singleAdd_a_6;
    _zz_singleAdd_a_8 <= _zz_singleAdd_a_7;
    _zz_singleAdd_a_9 <= _zz_singleAdd_a_8;
    _zz_singleAdd_a_10 <= _zz_singleAdd_a_9;
    _zz_singleAdd_a_11 <= io_a[191 : 128];
    _zz_singleAdd_a_12 <= _zz_singleAdd_a_11;
    _zz_singleAdd_a_13 <= _zz_singleAdd_a_12;
    _zz_singleAdd_a_14 <= _zz_singleAdd_a_13;
    _zz_singleAdd_a_15 <= io_a[255 : 192];
    _zz_singleAdd_a_16 <= _zz_singleAdd_a_15;
    _zz_singleAdd_a_17 <= _zz_singleAdd_a_16;
    _zz_singleAdd_a_18 <= io_a[319 : 256];
    _zz_singleAdd_a_19 <= _zz_singleAdd_a_18;
    _zz_singleAdd_a_20 <= io_a[377 : 320];
    _zz_io_r <= (singleAdd_add_io_s[377] ? _zz__zz_io_r : _zz__zz_io_r_1);
  end


endmodule

module BADD_9 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  input               io_c,
  output reg [377:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [64:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_5;
  wire       [64:0]   _zz__zz_io_s_5_1;
  wire       [0:0]    _zz__zz_io_s_5_2;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [64:0]   _zz__zz_io_s_32;
  wire       [64:0]   _zz__zz_io_s_32_1;
  wire       [0:0]    _zz__zz_io_s_32_2;
  wire       [57:0]   _zz__zz_io_s_45;
  wire       [57:0]   _zz__zz_io_s_45_1;
  wire       [0:0]    _zz__zz_io_s_45_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  wire       [64:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg        [63:0]   _zz_io_s_25;
  reg        [63:0]   _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg        [63:0]   _zz_io_s_29;
  reg        [63:0]   _zz_io_s_30;
  reg        [63:0]   _zz_io_s_31;
  wire       [64:0]   _zz_io_s_32;
  reg        [63:0]   _zz_io_s_33;
  reg                 _zz_io_s_34;
  reg        [56:0]   _zz_io_s_35;
  reg        [56:0]   _zz_io_s_36;
  reg        [56:0]   _zz_io_s_37;
  reg        [56:0]   _zz_io_s_38;
  reg        [56:0]   _zz_io_s_39;
  reg        [56:0]   _zz_io_s_40;
  reg        [56:0]   _zz_io_s_41;
  reg        [56:0]   _zz_io_s_42;
  reg        [56:0]   _zz_io_s_43;
  reg        [56:0]   _zz_io_s_44;
  wire       [57:0]   _zz_io_s_45;
  reg        [56:0]   _zz_io_s_46;
  reg                 _zz_io_s_47;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,io_b[63 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {64'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_5 = ({1'b0,_zz_io_s_3} + {1'b0,_zz_io_s_4});
  assign _zz__zz_io_s_5_2 = _zz_io_s_2;
  assign _zz__zz_io_s_5_1 = {64'd0, _zz__zz_io_s_5_2};
  assign _zz__zz_io_s_12 = ({1'b0,_zz_io_s_9} + {1'b0,_zz_io_s_11});
  assign _zz__zz_io_s_12_2 = _zz_io_s_7;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_17} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_14;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_32 = ({1'b0,_zz_io_s_27} + {1'b0,_zz_io_s_31});
  assign _zz__zz_io_s_32_2 = _zz_io_s_23;
  assign _zz__zz_io_s_32_1 = {64'd0, _zz__zz_io_s_32_2};
  assign _zz__zz_io_s_45 = ({1'b0,_zz_io_s_39} + {1'b0,_zz_io_s_44});
  assign _zz__zz_io_s_45_2 = _zz_io_s_34;
  assign _zz__zz_io_s_45_1 = {57'd0, _zz__zz_io_s_45_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_1;
    io_s[127 : 64] = _zz_io_s_6;
    io_s[191 : 128] = _zz_io_s_13;
    io_s[255 : 192] = _zz_io_s_22;
    io_s[319 : 256] = _zz_io_s_33;
    io_s[376 : 320] = _zz_io_s_46;
    io_s[377] = _zz_io_s_47;
  end

  assign _zz_io_s_5 = (_zz__zz_io_s_5 + _zz__zz_io_s_5_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_32 = (_zz__zz_io_s_32 + _zz__zz_io_s_32_1);
  assign _zz_io_s_45 = (_zz__zz_io_s_45 + _zz__zz_io_s_45_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s[64];
    _zz_io_s_3 <= io_a[127 : 64];
    _zz_io_s_4 <= io_b[127 : 64];
    _zz_io_s_6 <= _zz_io_s_5[63:0];
    _zz_io_s_7 <= _zz_io_s_5[64];
    _zz_io_s_8 <= io_a[191 : 128];
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= io_b[191 : 128];
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_15 <= io_a[255 : 192];
    _zz_io_s_16 <= _zz_io_s_15;
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= io_b[255 : 192];
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_21[64];
    _zz_io_s_24 <= io_a[319 : 256];
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_25;
    _zz_io_s_27 <= _zz_io_s_26;
    _zz_io_s_28 <= io_b[319 : 256];
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz_io_s_29;
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_33 <= _zz_io_s_32[63:0];
    _zz_io_s_34 <= _zz_io_s_32[64];
    _zz_io_s_35 <= io_a[376 : 320];
    _zz_io_s_36 <= _zz_io_s_35;
    _zz_io_s_37 <= _zz_io_s_36;
    _zz_io_s_38 <= _zz_io_s_37;
    _zz_io_s_39 <= _zz_io_s_38;
    _zz_io_s_40 <= io_b[376 : 320];
    _zz_io_s_41 <= _zz_io_s_40;
    _zz_io_s_42 <= _zz_io_s_41;
    _zz_io_s_43 <= _zz_io_s_42;
    _zz_io_s_44 <= _zz_io_s_43;
    _zz_io_s_46 <= _zz_io_s_45[56:0];
    _zz_io_s_47 <= _zz_io_s_45[57];
  end


endmodule

//FineReduction_9 replaced by FineReduction_17

//BADD_10 replaced by BADD_18

//BCMUL replaced by BCMUL_8

//KaratsubaMUL_1 replaced by KaratsubaMUL_17

//KaratsubaMUL replaced by KaratsubaMUL_16

//FineReduction_10 replaced by FineReduction_17

//BADD_11 replaced by BADD_18

//BCMUL_1 replaced by BCMUL_8

//KaratsubaMUL_3 replaced by KaratsubaMUL_17

//KaratsubaMUL_2 replaced by KaratsubaMUL_16

//FineReduction_11 replaced by FineReduction_17

//BADD_12 replaced by BADD_18

//BCMUL_2 replaced by BCMUL_8

//KaratsubaMUL_5 replaced by KaratsubaMUL_17

//KaratsubaMUL_4 replaced by KaratsubaMUL_16

//FineReduction_12 replaced by FineReduction_17

//BADD_13 replaced by BADD_18

//BCMUL_3 replaced by BCMUL_8

//KaratsubaMUL_7 replaced by KaratsubaMUL_17

//KaratsubaMUL_6 replaced by KaratsubaMUL_16

//FineReduction_13 replaced by FineReduction_17

//BADD_14 replaced by BADD_18

//BCMUL_4 replaced by BCMUL_8

//KaratsubaMUL_9 replaced by KaratsubaMUL_17

//KaratsubaMUL_8 replaced by KaratsubaMUL_16

//FineReduction_14 replaced by FineReduction_17

//BADD_15 replaced by BADD_18

//BCMUL_5 replaced by BCMUL_8

//KaratsubaMUL_11 replaced by KaratsubaMUL_17

//KaratsubaMUL_10 replaced by KaratsubaMUL_16

//FineReduction_15 replaced by FineReduction_17

//BADD_16 replaced by BADD_18

//BCMUL_6 replaced by BCMUL_8

//KaratsubaMUL_13 replaced by KaratsubaMUL_17

//KaratsubaMUL_12 replaced by KaratsubaMUL_16

//FineReduction_16 replaced by FineReduction_17

//BADD_17 replaced by BADD_18

//BCMUL_7 replaced by BCMUL_8

//KaratsubaMUL_15 replaced by KaratsubaMUL_17

//KaratsubaMUL_14 replaced by KaratsubaMUL_16

module FineReduction_17 (
  input      [378:0]  io_a,
  output     [376:0]  io_r,
  input               clk,
  input               resetn
);

  wire       [377:0]  doubleAdd_reduction_io_a;
  wire       [378:0]  doubleAdd_add_io_s;
  wire       [376:0]  doubleAdd_reduction_io_r;
  wire       [376:0]  _zz_doubleAdd_subRom_1;
  wire       [376:0]  _zz_doubleAdd_subRom_2;
  wire       [377:0]  _zz_doubleAdd_subRom_3;
  wire       [377:0]  _zz_doubleAdd_subRom_4;
  wire       [376:0]  _zz_doubleAdd_subRom_5;
  reg        [377:0]  _zz__zz_io_b;
  wire       [2:0]    _zz__zz_io_b_1;
  wire       [377:0]  doubleAdd_subRom_0;
  wire       [377:0]  doubleAdd_subRom_1;
  wire       [377:0]  doubleAdd_subRom_2;
  wire       [377:0]  doubleAdd_subRom_3;
  wire       [377:0]  doubleAdd_subRom_4;
  wire       [377:0]  doubleAdd_subRom_5;
  wire       [377:0]  doubleAdd_subRom_6;
  wire       [377:0]  doubleAdd_subRom_7;
  reg        [377:0]  _zz_io_a;
  reg        [377:0]  _zz_io_b;

  assign _zz_doubleAdd_subRom_1 = 377'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001;
  assign _zz_doubleAdd_subRom_2 = 377'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001;
  assign _zz_doubleAdd_subRom_3 = 378'h35c748c2f8a21d58c760b80d94292763445b3e601ea271e3de6c45f741290002e16ba88600000010a11800000000002;
  assign _zz_doubleAdd_subRom_4 = 378'h35c748c2f8a21d58c760b80d94292763445b3e601ea271e3de6c45f741290002e16ba88600000010a11800000000002;
  assign _zz_doubleAdd_subRom_5 = 377'h10aaed2474f32c052b1114145e3dbb14e688dd902df3aad5cda268f2e1bd800452217cc900000018f1a400000000003;
  assign _zz__zz_io_b_1 = io_a[378 : 376];
  BADD_531 doubleAdd_add (
    .io_a   (_zz_io_a[377:0]          ), //i
    .io_b   (_zz_io_b[377:0]          ), //i
    .io_c   (1'b1                     ), //i
    .io_s   (doubleAdd_add_io_s[378:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  FineReduction_26 doubleAdd_reduction (
    .io_a   (doubleAdd_reduction_io_a[377:0]), //i
    .io_r   (doubleAdd_reduction_io_r[376:0]), //o
    .clk    (clk                            ), //i
    .resetn (resetn                         )  //i
  );
  always @(*) begin
    case(_zz__zz_io_b_1)
      3'b000 : _zz__zz_io_b = doubleAdd_subRom_0;
      3'b001 : _zz__zz_io_b = doubleAdd_subRom_1;
      3'b010 : _zz__zz_io_b = doubleAdd_subRom_2;
      3'b011 : _zz__zz_io_b = doubleAdd_subRom_3;
      3'b100 : _zz__zz_io_b = doubleAdd_subRom_4;
      3'b101 : _zz__zz_io_b = doubleAdd_subRom_5;
      3'b110 : _zz__zz_io_b = doubleAdd_subRom_6;
      default : _zz__zz_io_b = doubleAdd_subRom_7;
    endcase
  end

  assign doubleAdd_subRom_0 = 378'h0;
  assign doubleAdd_subRom_1 = {1'd0, _zz_doubleAdd_subRom_1};
  assign doubleAdd_subRom_2 = {1'd0, _zz_doubleAdd_subRom_2};
  assign doubleAdd_subRom_3 = _zz_doubleAdd_subRom_3;
  assign doubleAdd_subRom_4 = _zz_doubleAdd_subRom_4;
  assign doubleAdd_subRom_5 = {1'd0, _zz_doubleAdd_subRom_5};
  assign doubleAdd_subRom_6 = 378'h0;
  assign doubleAdd_subRom_7 = 378'h0;
  assign doubleAdd_reduction_io_a = doubleAdd_add_io_s[377:0];
  assign io_r = doubleAdd_reduction_io_r;
  always @(posedge clk) begin
    _zz_io_a <= io_a[377:0];
    _zz_io_b <= _zz__zz_io_b;
  end


endmodule

module BADD_18 (
  input      [378:0]  io_a,
  input      [378:0]  io_b,
  input               io_c,
  output reg [379:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [378:0]  _zz__zz_io_s_1;
  wire       [64:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [378:0]  _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_10;
  wire       [64:0]   _zz__zz_io_s_10_1;
  wire       [0:0]    _zz__zz_io_s_10_2;
  wire       [378:0]  _zz__zz_io_s_19;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [378:0]  _zz__zz_io_s_30;
  wire       [64:0]   _zz__zz_io_s_33;
  wire       [64:0]   _zz__zz_io_s_33_1;
  wire       [0:0]    _zz__zz_io_s_33_2;
  wire       [378:0]  _zz__zz_io_s_42;
  wire       [64:0]   _zz__zz_io_s_46;
  wire       [64:0]   _zz__zz_io_s_46_1;
  wire       [0:0]    _zz__zz_io_s_46_2;
  wire       [378:0]  _zz__zz_io_s_55;
  wire       [59:0]   _zz__zz_io_s_60;
  wire       [59:0]   _zz__zz_io_s_60_1;
  wire       [0:0]    _zz__zz_io_s_60_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  wire       [64:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg        [63:0]   _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg                 _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg        [63:0]   _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg        [63:0]   _zz_io_s_25;
  reg                 _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg        [63:0]   _zz_io_s_29;
  reg        [63:0]   _zz_io_s_30;
  reg        [63:0]   _zz_io_s_31;
  reg        [63:0]   _zz_io_s_32;
  wire       [64:0]   _zz_io_s_33;
  reg        [63:0]   _zz_io_s_34;
  reg        [63:0]   _zz_io_s_35;
  reg        [63:0]   _zz_io_s_36;
  reg                 _zz_io_s_37;
  reg        [63:0]   _zz_io_s_38;
  reg        [63:0]   _zz_io_s_39;
  reg        [63:0]   _zz_io_s_40;
  reg        [63:0]   _zz_io_s_41;
  reg        [63:0]   _zz_io_s_42;
  reg        [63:0]   _zz_io_s_43;
  reg        [63:0]   _zz_io_s_44;
  reg        [63:0]   _zz_io_s_45;
  wire       [64:0]   _zz_io_s_46;
  reg        [63:0]   _zz_io_s_47;
  reg        [63:0]   _zz_io_s_48;
  reg                 _zz_io_s_49;
  reg        [58:0]   _zz_io_s_50;
  reg        [58:0]   _zz_io_s_51;
  reg        [58:0]   _zz_io_s_52;
  reg        [58:0]   _zz_io_s_53;
  reg        [58:0]   _zz_io_s_54;
  reg        [58:0]   _zz_io_s_55;
  reg        [58:0]   _zz_io_s_56;
  reg        [58:0]   _zz_io_s_57;
  reg        [58:0]   _zz_io_s_58;
  reg        [58:0]   _zz_io_s_59;
  wire       [59:0]   _zz_io_s_60;
  reg        [58:0]   _zz_io_s_61;
  reg                 _zz_io_s_62;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,_zz__zz_io_s_1[63 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {64'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_9 = (~ io_b);
  assign _zz__zz_io_s_10 = ({1'b0,_zz_io_s_8} + {1'b0,_zz_io_s_9});
  assign _zz__zz_io_s_10_2 = _zz_io_s_7;
  assign _zz__zz_io_s_10_1 = {64'd0, _zz__zz_io_s_10_2};
  assign _zz__zz_io_s_19 = (~ io_b);
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_18} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_16;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_30 = (~ io_b);
  assign _zz__zz_io_s_33 = ({1'b0,_zz_io_s_29} + {1'b0,_zz_io_s_32});
  assign _zz__zz_io_s_33_2 = _zz_io_s_26;
  assign _zz__zz_io_s_33_1 = {64'd0, _zz__zz_io_s_33_2};
  assign _zz__zz_io_s_42 = (~ io_b);
  assign _zz__zz_io_s_46 = ({1'b0,_zz_io_s_41} + {1'b0,_zz_io_s_45});
  assign _zz__zz_io_s_46_2 = _zz_io_s_37;
  assign _zz__zz_io_s_46_1 = {64'd0, _zz__zz_io_s_46_2};
  assign _zz__zz_io_s_55 = (~ io_b);
  assign _zz__zz_io_s_60 = ({1'b0,_zz_io_s_54} + {1'b0,_zz_io_s_59});
  assign _zz__zz_io_s_60_2 = _zz_io_s_49;
  assign _zz__zz_io_s_60_1 = {59'd0, _zz__zz_io_s_60_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_6;
    io_s[127 : 64] = _zz_io_s_15;
    io_s[191 : 128] = _zz_io_s_25;
    io_s[255 : 192] = _zz_io_s_36;
    io_s[319 : 256] = _zz_io_s_48;
    io_s[378 : 320] = _zz_io_s_61;
    io_s[379] = (! _zz_io_s_62);
  end

  assign _zz_io_s_10 = (_zz__zz_io_s_10 + _zz__zz_io_s_10_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_33 = (_zz__zz_io_s_33 + _zz__zz_io_s_33_1);
  assign _zz_io_s_46 = (_zz__zz_io_s_46 + _zz__zz_io_s_46_1);
  assign _zz_io_s_60 = (_zz__zz_io_s_60 + _zz__zz_io_s_60_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= _zz_io_s[64];
    _zz_io_s_8 <= io_a[127 : 64];
    _zz_io_s_9 <= _zz__zz_io_s_9[127 : 64];
    _zz_io_s_11 <= _zz_io_s_10[63:0];
    _zz_io_s_12 <= _zz_io_s_11;
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_13;
    _zz_io_s_15 <= _zz_io_s_14;
    _zz_io_s_16 <= _zz_io_s_10[64];
    _zz_io_s_17 <= io_a[191 : 128];
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= _zz__zz_io_s_19[191 : 128];
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_22;
    _zz_io_s_24 <= _zz_io_s_23;
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_21[64];
    _zz_io_s_27 <= io_a[255 : 192];
    _zz_io_s_28 <= _zz_io_s_27;
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz__zz_io_s_30[255 : 192];
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_32 <= _zz_io_s_31;
    _zz_io_s_34 <= _zz_io_s_33[63:0];
    _zz_io_s_35 <= _zz_io_s_34;
    _zz_io_s_36 <= _zz_io_s_35;
    _zz_io_s_37 <= _zz_io_s_33[64];
    _zz_io_s_38 <= io_a[319 : 256];
    _zz_io_s_39 <= _zz_io_s_38;
    _zz_io_s_40 <= _zz_io_s_39;
    _zz_io_s_41 <= _zz_io_s_40;
    _zz_io_s_42 <= _zz__zz_io_s_42[319 : 256];
    _zz_io_s_43 <= _zz_io_s_42;
    _zz_io_s_44 <= _zz_io_s_43;
    _zz_io_s_45 <= _zz_io_s_44;
    _zz_io_s_47 <= _zz_io_s_46[63:0];
    _zz_io_s_48 <= _zz_io_s_47;
    _zz_io_s_49 <= _zz_io_s_46[64];
    _zz_io_s_50 <= io_a[378 : 320];
    _zz_io_s_51 <= _zz_io_s_50;
    _zz_io_s_52 <= _zz_io_s_51;
    _zz_io_s_53 <= _zz_io_s_52;
    _zz_io_s_54 <= _zz_io_s_53;
    _zz_io_s_55 <= _zz__zz_io_s_55[378 : 320];
    _zz_io_s_56 <= _zz_io_s_55;
    _zz_io_s_57 <= _zz_io_s_56;
    _zz_io_s_58 <= _zz_io_s_57;
    _zz_io_s_59 <= _zz_io_s_58;
    _zz_io_s_61 <= _zz_io_s_60[58:0];
    _zz_io_s_62 <= _zz_io_s_60[59];
  end


endmodule

module BCMUL_8 (
  input      [377:0]  io_a,
  output     [378:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [322:0]  NAFElements_adds_0_io_a;
  wire       [322:0]  NAFElements_adds_0_io_b;
  wire       [332:0]  NAFElements_adds_1_io_a;
  wire       [332:0]  NAFElements_adds_1_io_b;
  wire       [272:0]  NAFElements_adds_2_io_a;
  wire       [272:0]  NAFElements_adds_2_io_b;
  wire       [189:0]  NAFElements_adds_3_io_a;
  wire       [189:0]  NAFElements_adds_3_io_b;
  wire       [327:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [280:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [315:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [253:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [234:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [209:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [170:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [176:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [214:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [116:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [136:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [106:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [91:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [101:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [111:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [50:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [25:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [15:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [20:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [31:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [4:0]    adder_posMUL_multiElements_add_add_io_a;
  wire       [267:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [225:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [258:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [194:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [200:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [220:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [182:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [150:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [166:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [141:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [125:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [129:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [145:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [74:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [84:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [63:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [54:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [58:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [68:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a;
  wire       [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_a;
  wire       [120:0]  adder_negMUL_multiElements_add_add_io_a;
  wire       [378:0]  adder_add_io_b;
  wire       [323:0]  NAFElements_adds_0_io_s;
  wire       [333:0]  NAFElements_adds_1_io_s;
  wire       [273:0]  NAFElements_adds_2_io_s;
  wire       [190:0]  NAFElements_adds_3_io_s;
  wire       [333:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [323:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [328:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [287:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [277:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [281:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [316:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [254:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [235:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [240:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [210:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [171:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [177:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [215:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [263:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [155:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [117:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [137:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [107:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [92:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [102:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [112:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [51:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [43:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [47:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [26:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [16:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [21:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [32:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [80:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [163:0]  adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [5:0]    adder_posMUL_multiElements_add_add_io_s;
  wire       [268:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [226:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [259:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [206:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [195:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [201:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [221:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [183:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [151:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [167:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [142:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [126:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [130:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [146:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [190:0]  adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [97:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [75:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [85:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [64:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [55:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [59:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [69:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s;
  wire       [10:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [37:0]   adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_s;
  wire       [121:0]  adder_negMUL_multiElements_add_add_io_s;
  wire       [379:0]  adder_add_io_s;
  wire       [379:0]  _zz_io_a_11;
  wire       [378:0]  _zz_io_a_12;
  wire       [380:0]  _zz_io_a_13;
  wire       [380:0]  _zz_io_a_14;
  wire       [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  wire       [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  wire       [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  wire       [12:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  wire       [12:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  wire       [12:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  wire       [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  wire       [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  wire       [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  wire       [0:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  wire       [0:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  wire       [0:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  wire       [50:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [46:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [42:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [31:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [25:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [20:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [15:0]   _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [4:0]    _zz__zz_adder_posMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [58:0]   _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [54:0]   _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [36:0]   _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [9:0]    _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [378:0]  _zz_io_p;
  wire       [379:0]  _zz_io_p_1;
  wire       [378:0]  _zz_NAFElements_sums_0;
  reg        [63:0]   _zz_NAFElements_sums_0_1;
  reg        [63:0]   _zz_NAFElements_sums_0_2;
  reg        [63:0]   _zz_NAFElements_sums_0_3;
  reg        [63:0]   _zz_NAFElements_sums_0_4;
  reg        [63:0]   _zz_NAFElements_sums_0_5;
  reg        [63:0]   _zz_NAFElements_sums_0_6;
  reg        [63:0]   _zz_NAFElements_sums_0_7;
  reg        [63:0]   _zz_NAFElements_sums_0_8;
  reg        [63:0]   _zz_NAFElements_sums_0_9;
  reg        [63:0]   _zz_NAFElements_sums_0_10;
  reg        [58:0]   _zz_NAFElements_sums_0_11;
  reg        [58:0]   _zz_NAFElements_sums_0_12;
  reg        [58:0]   _zz_NAFElements_sums_0_13;
  reg        [58:0]   _zz_NAFElements_sums_0_14;
  reg        [58:0]   _zz_NAFElements_sums_0_15;
  wire       [378:0]  NAFElements_sums_0;
  wire       [322:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [332:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [272:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [189:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [378:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [378:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [332:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [332:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [332:0]  _zz_io_a;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [45:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [327:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [327:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [327:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  wire       [322:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [322:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [55:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [322:0]  _zz_io_a_1;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [315:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [315:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [315:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [315:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  wire       [59:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [58:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  wire       [286:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [286:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [286:0]  _zz_io_a_2;
  reg        [28:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [28:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [280:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [280:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [280:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [29:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [29:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [29:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [33:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [29:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [24:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  wire       [276:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [276:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [276:0]  _zz_io_a_3;
  reg        [3:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [3:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [34:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [62:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [262:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [262:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [11:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [11:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [11:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [51:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [11:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [6:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  wire       [253:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [253:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  wire       [61:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [2:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [2:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [60:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [2:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [58:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [58:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [2:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [8:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [239:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [239:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [239:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20;
  wire       [234:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [234:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [239:0]  _zz_io_a_4;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [214:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [214:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [214:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [214:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [35:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20;
  wire       [209:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [209:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [40:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [22:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [17:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20;
  reg        [209:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [176:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [176:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [176:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [53:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [48:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [48:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [48:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  wire       [170:0]  adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [170:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [115:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [162:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [162:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [23:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [39:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [34:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [34:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [34:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  wire       [154:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [154:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [26:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [26:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [26:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [154:0]  _zz_io_a_5;
  reg        [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [7:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [136:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [136:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [136:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [49:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [13:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [8:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [8:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [8:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  wire       [116:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [116:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [57:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [57:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [57:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [57:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [19:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [111:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [111:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [111:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [111:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [52:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  wire       [106:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [106:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [106:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [101:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [101:0]  adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [101:0]  _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [37:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  wire       [91:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [91:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [30:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [27:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [91:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [9:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [79:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [79:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  wire       [50:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [50:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [28:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [46:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [46:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [46:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [42:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [42:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [42:0]   _zz_io_a_6;
  reg        [3:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [3:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [46:0]   _zz_io_a_7;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [32:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [31:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [31:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [31:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [31:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  wire       [25:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [25:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [5:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [20:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [20:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [20:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [15:0]   adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [15:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [4:0]    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [10:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [47:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [82:0]   _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [215:0]  _zz_adder_posMUL_multiElements_lsbMUL_p;
  wire       [4:0]    adder_posMUL_multiElements_msbMUL_p;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p_1;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p_2;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p_3;
  reg        [4:0]    _zz_adder_posMUL_multiElements_msbMUL_p_4;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_1;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_2;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_3;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_4;
  reg        [4:0]    adder_posMUL_multiElements_msbMUL_p_delay_5;
  reg        [373:0]  _zz_adder_posMUL_p;
  reg        [272:0]  adder_negMUL_p;
  reg        [272:0]  adder_negMUL_multiElements_lsbMUL_p;
  reg        [272:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [272:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [272:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [272:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [272:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [21:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [21:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [21:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [41:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [21:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  wire       [267:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [267:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [46:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [16:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [11:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [4:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [258:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [258:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [258:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  wire       [225:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [225:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [24:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20;
  reg        [32:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [220:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [220:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [220:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [220:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [29:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [33:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [28:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  reg        [28:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20;
  wire       [205:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [205:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20;
  reg        [205:0]  _zz_io_a_8;
  reg        [14:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [14:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [200:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [200:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [200:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [49:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [8:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  reg        [8:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20;
  wire       [194:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [194:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [55:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [7:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20;
  reg        [194:0]  adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
  reg        [5:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [51:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [189:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [189:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  wire       [61:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  wire       [182:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [182:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [59:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [54:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [54:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [54:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [166:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [166:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [166:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [19:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [38:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  wire       [150:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [150:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [35:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [27:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
  reg        [15:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [166:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [145:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [145:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [145:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [145:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [40:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
  reg        [22:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
  reg        [17:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
  reg        [17:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
  reg        [17:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
  wire       [141:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [141:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [44:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
  reg        [18:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
  reg        [13:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [129:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [129:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [129:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [56:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
  reg        [6:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16;
  reg        [1:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
  reg        [1:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
  reg        [1:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
  wire       [125:0]  adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [125:0]  _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  wire       [61:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [60:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [58:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
  reg        [2:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16;
  reg        [3:0]    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [15:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [43:0]   _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [82:0]   _zz_adder_negMUL_multiElements_lsbMUL_p;
  reg        [120:0]  adder_negMUL_multiElements_msbMUL_p;
  reg        [120:0]  adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [120:0]  adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [120:0]  adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [120:0]  adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [120:0]  _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [1:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [61:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [61:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [61:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [61:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [56:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [56:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [56:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [56:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  wire       [96:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [96:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
  reg        [32:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
  reg        [32:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
  reg        [32:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
  reg        [32:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
  reg        [96:0]   _zz_io_a_9;
  reg        [23:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [23:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [84:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [84:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [84:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
  reg        [37:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
  reg        [25:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
  reg        [20:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
  reg        [20:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
  reg        [20:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
  reg        [20:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
  wire       [74:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [74:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
  reg        [47:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6;
  reg        [15:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
  reg        [15:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
  reg        [15:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
  reg        [15:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
  reg        [10:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
  reg        [10:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
  reg        [10:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
  reg        [10:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [35:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  reg        [68:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [68:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  wire       [68:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [68:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
  reg        [53:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
  wire       [63:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  wire       [63:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
  reg        [4:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [58:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [58:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [58:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [54:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [54:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [54:0]   adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
  reg        [3:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  reg        [51:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  wire       [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
  reg        [36:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  wire       [9:0]    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
  reg        [9:0]    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  reg        [9:0]    _zz_io_a_10;
  reg        [26:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  reg        [26:0]   _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
  reg        [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
  reg        [36:0]   adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_2;
  reg        [83:0]   _zz_adder_negMUL_multiElements_msbMUL_p;
  reg        [151:0]  _zz_adder_negMUL_p;
  reg        [272:0]  adder_negMUL_p_delay_1;

  assign _zz_io_a_11 = ({2'd0,io_a} <<< 2);
  assign _zz_io_a_12 = ({1'd0,io_a} <<< 1);
  assign _zz_io_a_13 = ({3'd0,io_a} <<< 3);
  assign _zz_io_a_14 = ({3'd0,io_a} <<< 3);
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_sums_0[50:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[46:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[42:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[31:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[25:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[20:0];
  assign _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[15:0];
  assign _zz__zz_adder_posMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[58:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_sums_0[54:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[36:0];
  assign _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[9:0];
  assign _zz_io_p_1 = adder_add_io_s;
  assign _zz_io_p = _zz_io_p_1[378:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[17 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[17 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[17 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[12 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[12 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[12 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4[7 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[7 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[7 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[0 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[0 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[0 : 0];
  BADD_532 NAFElements_adds_0 (
    .io_a   (NAFElements_adds_0_io_a[322:0]), //i
    .io_b   (NAFElements_adds_0_io_b[322:0]), //i
    .io_c   (1'b0                          ), //i
    .io_s   (NAFElements_adds_0_io_s[323:0]), //o
    .clk    (clk                           ), //i
    .resetn (resetn                        )  //i
  );
  BADD_533 NAFElements_adds_1 (
    .io_a   (NAFElements_adds_1_io_a[332:0]), //i
    .io_b   (NAFElements_adds_1_io_b[332:0]), //i
    .io_c   (1'b0                          ), //i
    .io_s   (NAFElements_adds_1_io_s[333:0]), //o
    .clk    (clk                           ), //i
    .resetn (resetn                        )  //i
  );
  BADD_534 NAFElements_adds_2 (
    .io_a   (NAFElements_adds_2_io_a[272:0]), //i
    .io_b   (NAFElements_adds_2_io_b[272:0]), //i
    .io_c   (1'b0                          ), //i
    .io_s   (NAFElements_adds_2_io_s[273:0]), //o
    .clk    (clk                           ), //i
    .resetn (resetn                        )  //i
  );
  BADD_535 NAFElements_adds_3 (
    .io_a   (NAFElements_adds_3_io_a[189:0]), //i
    .io_b   (NAFElements_adds_3_io_b[189:0]), //i
    .io_c   (1'b1                          ), //i
    .io_s   (NAFElements_adds_3_io_s[190:0]), //o
    .clk    (clk                           ), //i
    .resetn (resetn                        )  //i
  );
  BADD_536 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a[332:0]                                                                                                                                        ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[332:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[333:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_537 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_1[322:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[322:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[323:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_538 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[327:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[327:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[328:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_539 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_2[286:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[286:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[287:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_540 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_3[276:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[276:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[277:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_541 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[280:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[280:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[281:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_542 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[315:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[315:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[316:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_543 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[253:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[253:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[254:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_544 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[234:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[234:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[235:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_545 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_4[239:0]                                                                                                                 ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[239:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[240:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_546 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[209:0]    ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1[209:0]), //i
    .io_c   (1'b0                                                                                                                                                       ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[210:0]    ), //o
    .clk    (clk                                                                                                                                                        ), //i
    .resetn (resetn                                                                                                                                                     )  //i
  );
  BADD_547 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[170:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[170:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[171:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_548 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[176:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[176:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[177:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_549 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[214:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[214:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[215:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_550 adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[262:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[262:0]    ), //i
    .io_c   (1'b0                                                                                    ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[263:0]), //o
    .clk    (clk                                                                                     ), //i
    .resetn (resetn                                                                                  )  //i
  );
  BADD_551 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_5[154:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[154:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[155:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_552 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[116:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[116:0]    ), //i
    .io_c   (1'b0                                                                                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[117:0]), //o
    .clk    (clk                                                                                                                                                    ), //i
    .resetn (resetn                                                                                                                                                 )  //i
  );
  BADD_553 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[136:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[136:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[137:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_554 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[106:0]    ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1[106:0]), //i
    .io_c   (1'b0                                                                                                                                                       ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[107:0]    ), //o
    .clk    (clk                                                                                                                                                        ), //i
    .resetn (resetn                                                                                                                                                     )  //i
  );
  BADD_555 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[91:0]    ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1[91:0]), //i
    .io_c   (1'b0                                                                                                                                                      ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[92:0]    ), //o
    .clk    (clk                                                                                                                                                       ), //i
    .resetn (resetn                                                                                                                                                    )  //i
  );
  BADD_556 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[101:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[101:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[102:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_557 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[111:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[111:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[112:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_558 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[50:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[50:0]    ), //i
    .io_c   (1'b0                                                                                                                                                  ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[51:0]), //o
    .clk    (clk                                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                                )  //i
  );
  BADD_559 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_6[42:0]                                                                                                                                      ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[42:0]    ), //i
    .io_c   (1'b0                                                                                                                                                  ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[43:0]), //o
    .clk    (clk                                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                                )  //i
  );
  BADD_560 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_7[46:0]                                                                                                                 ), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[46:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[47:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_561 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[25:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[25:0]    ), //i
    .io_c   (1'b0                                                                                                                                                  ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[26:0]), //o
    .clk    (clk                                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                                )  //i
  );
  BADD_562 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[15:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[15:0]    ), //i
    .io_c   (1'b0                                                                                                                                                  ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[16:0]), //o
    .clk    (clk                                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                                )  //i
  );
  BADD_563 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[20:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[20:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[21:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_564 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[31:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[31:0]    ), //i
    .io_c   (1'b0                                                                                                        ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[32:0]), //o
    .clk    (clk                                                                                                         ), //i
    .resetn (resetn                                                                                                      )  //i
  );
  BADD_565 adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[79:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[79:0]    ), //i
    .io_c   (1'b0                                                                                   ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[80:0]), //o
    .clk    (clk                                                                                    ), //i
    .resetn (resetn                                                                                 )  //i
  );
  BADD_566 adder_posMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_a[162:0]), //i
    .io_b   (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p[162:0]    ), //i
    .io_c   (1'b0                                                               ), //i
    .io_s   (adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_s[163:0]), //o
    .clk    (clk                                                                ), //i
    .resetn (resetn                                                             )  //i
  );
  BADD_567 adder_posMUL_multiElements_add_add (
    .io_a   (adder_posMUL_multiElements_add_add_io_a[4:0]    ), //i
    .io_b   (adder_posMUL_multiElements_msbMUL_p_delay_5[4:0]), //i
    .io_c   (1'b0                                            ), //i
    .io_s   (adder_posMUL_multiElements_add_add_io_s[5:0]    ), //o
    .clk    (clk                                             ), //i
    .resetn (resetn                                          )  //i
  );
  BADD_568 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[267:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[267:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[268:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_569 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[225:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[225:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[226:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_570 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[258:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[258:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[259:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_571 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_8[205:0]                                                                                                                 ), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[205:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[206:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_572 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[194:0]    ), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1[194:0]), //i
    .io_c   (1'b0                                                                                                                                  ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[195:0]    ), //o
    .clk    (clk                                                                                                                                   ), //i
    .resetn (resetn                                                                                                                                )  //i
  );
  BADD_573 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[200:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[200:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[201:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_574 adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[220:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[220:0]    ), //i
    .io_c   (1'b0                                                                                    ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[221:0]), //o
    .clk    (clk                                                                                     ), //i
    .resetn (resetn                                                                                  )  //i
  );
  BADD_575 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[182:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[182:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[183:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_576 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[150:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[150:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[151:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_577 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[166:0]    ), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1[166:0]), //i
    .io_c   (1'b0                                                                                                             ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[167:0]    ), //o
    .clk    (clk                                                                                                              ), //i
    .resetn (resetn                                                                                                           )  //i
  );
  BADD_578 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[141:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[141:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[142:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_579 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[125:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[125:0]    ), //i
    .io_c   (1'b0                                                                                                                              ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[126:0]), //o
    .clk    (clk                                                                                                                               ), //i
    .resetn (resetn                                                                                                                            )  //i
  );
  BADD_580 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[129:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[129:0]    ), //i
    .io_c   (1'b0                                                                                                         ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[130:0]), //o
    .clk    (clk                                                                                                          ), //i
    .resetn (resetn                                                                                                       )  //i
  );
  BADD_581 adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[145:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[145:0]    ), //i
    .io_c   (1'b0                                                                                    ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[146:0]), //o
    .clk    (clk                                                                                     ), //i
    .resetn (resetn                                                                                  )  //i
  );
  BADD_582 adder_negMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_a[189:0]), //i
    .io_b   (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p[189:0]    ), //i
    .io_c   (1'b0                                                               ), //i
    .io_s   (adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_s[190:0]), //o
    .clk    (clk                                                                ), //i
    .resetn (resetn                                                             )  //i
  );
  BADD_583 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_9[96:0]                                                                                                                 ), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[96:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[97:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_584 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[74:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[74:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[75:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_585 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[84:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[84:0]    ), //i
    .io_c   (1'b0                                                                                                        ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[85:0]), //o
    .clk    (clk                                                                                                         ), //i
    .resetn (resetn                                                                                                      )  //i
  );
  BADD_586 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[63:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63:0]    ), //i
    .io_c   (1'b0                                                                                                                             ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[64:0]), //o
    .clk    (clk                                                                                                                              ), //i
    .resetn (resetn                                                                                                                           )  //i
  );
  BADD_587 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a[54:0]    ), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1[54:0]), //i
    .io_c   (1'b0                                                                                                                                 ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[55:0]    ), //o
    .clk    (clk                                                                                                                                  ), //i
    .resetn (resetn                                                                                                                               )  //i
  );
  BADD_588 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a[58:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[58:0]    ), //i
    .io_c   (1'b0                                                                                                        ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[59:0]), //o
    .clk    (clk                                                                                                         ), //i
    .resetn (resetn                                                                                                      )  //i
  );
  BADD_589 adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a[68:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[68:0]    ), //i
    .io_c   (1'b0                                                                                   ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[69:0]), //o
    .clk    (clk                                                                                    ), //i
    .resetn (resetn                                                                                 )  //i
  );
  BADD_590 adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (_zz_io_a_10[9:0]                                                                       ), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[9:0]     ), //i
    .io_c   (1'b0                                                                                   ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[10:0]), //o
    .clk    (clk                                                                                    ), //i
    .resetn (resetn                                                                                 )  //i
  );
  BADD_591 adder_negMUL_multiElements_msbMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_a[36:0]    ), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_2[36:0]), //i
    .io_c   (1'b0                                                                  ), //i
    .io_s   (adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_s[37:0]    ), //o
    .clk    (clk                                                                   ), //i
    .resetn (resetn                                                                )  //i
  );
  BADD_592 adder_negMUL_multiElements_add_add (
    .io_a   (adder_negMUL_multiElements_add_add_io_a[120:0]), //i
    .io_b   (adder_negMUL_multiElements_msbMUL_p[120:0]    ), //i
    .io_c   (1'b0                                          ), //i
    .io_s   (adder_negMUL_multiElements_add_add_io_s[121:0]), //o
    .clk    (clk                                           ), //i
    .resetn (resetn                                        )  //i
  );
  BADD_593 adder_add (
    .io_a   (adder_posMUL_p[378:0]), //i
    .io_b   (adder_add_io_b[378:0]), //i
    .io_c   (1'b1                 ), //i
    .io_s   (adder_add_io_s[379:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign NAFElements_adds_0_io_a = _zz_io_a_11[322:0];
  assign NAFElements_adds_0_io_b = io_a[322:0];
  assign NAFElements_adds_1_io_a = _zz_io_a_12[332:0];
  assign NAFElements_adds_1_io_b = io_a[332:0];
  assign NAFElements_adds_2_io_a = _zz_io_a_13[272:0];
  assign NAFElements_adds_2_io_b = io_a[272:0];
  assign NAFElements_adds_3_io_a = _zz_io_a_14[189:0];
  assign NAFElements_adds_3_io_b = io_a[189:0];
  assign _zz_NAFElements_sums_0 = {1'd0, io_a};
  assign NAFElements_sums_0 = {_zz_NAFElements_sums_0_15,{_zz_NAFElements_sums_0_10,{_zz_NAFElements_sums_0_6,{_zz_NAFElements_sums_0_3,{_zz_NAFElements_sums_0_1,_zz_NAFElements_sums_0[63 : 0]}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_adds_0_io_s[322:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_adds_1_io_s[332:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_adds_2_io_s[272:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_adds_3_io_s[189:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 320],{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[319 : 256],{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[255 : 192],{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128],{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64],_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0]}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[255 : 192];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[319 : 256];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[332 : 320],{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6[17 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5[17 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14}}}}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[45 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 46] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[332:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[327:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[255 : 192];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[319 : 256];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[327 : 320],{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5[12 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[12 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13}}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[255 : 192];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[319 : 256];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[322 : 320],{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6[7 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5[7 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14}}}}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[327 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[322:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 51);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[50 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 51] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[327:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[315:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[255 : 192];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[315 : 256];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5[0 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[0 : 0]},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[286:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[255 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7}}}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[28 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[315 : 29] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[286:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[280:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[255 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[276:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[255 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7}}}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[3 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[280 : 4] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[276:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 35);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[34 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[315 : 35] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[280:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 63);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[62 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 63] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[315:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[262:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[255 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7}}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_sums_0[253:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[253 : 192];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7}}}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 9);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[8 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[262 : 9] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[253:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[239:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[234:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8}}}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[239 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[234:0];
  end

  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[22 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[262 : 23] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[239:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[214:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8}}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_sums_0[209:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18},{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8}}}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[214 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[209:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[176:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[170:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9}}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 6);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[5 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[176 : 6] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[170:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 38);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[37 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[214 : 38] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[176:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 48);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[47 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[262 : 48] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[214:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 116);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[115 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[378 : 116] = adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[262:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[162:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[154:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9}}};
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[7 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[162 : 8] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[154:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[136:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[116:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 20);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[19 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[136 : 20] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[116:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 26);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[25 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[162 : 26] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[136:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[111:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = NAFElements_sums_0[106:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[111 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[106:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[101:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_sums_0[91:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 10);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[9 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[101 : 10] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[91:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 10);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[9 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[111 : 10] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[101:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 51);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[50 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[162 : 51] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[111:0];
  end

  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[79:0];
  assign _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14,{_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10}};
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 29);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[28 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[79 : 29] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[50:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[3 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[46 : 4] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[42:0];
  end

  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[32 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[79 : 33] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[46:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 6);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[5 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[31 : 6] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[25:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[4 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[20 : 5] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[15:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 11);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[10 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[31 : 11] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[20:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 48);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[47 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[79 : 48] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[31:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 83);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p[82 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p[162 : 83] = adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[79:0];
  end

  assign adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 216);
  always @(*) begin
    adder_posMUL_multiElements_lsbMUL_p[215 : 0] = _zz_adder_posMUL_multiElements_lsbMUL_p;
    adder_posMUL_multiElements_lsbMUL_p[378 : 216] = adder_posMUL_multiElements_lsbMUL_multiElements_add_add_io_s[162:0];
  end

  assign adder_posMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_msbMUL_p_4;
  assign adder_posMUL_multiElements_add_add_io_a = (adder_posMUL_multiElements_lsbMUL_p >>> 374);
  always @(*) begin
    adder_posMUL_p[373 : 0] = _zz_adder_posMUL_p;
    adder_posMUL_p[378 : 374] = adder_posMUL_multiElements_add_add_io_s[4:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[191 : 128];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[255 : 192];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8}}}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[267:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[255 : 192];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7}}}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[272 : 5] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[267:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[258:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[255 : 192];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7}}}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[225:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8}}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 33);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[32 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[258 : 33] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[225:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 14);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[13 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[272 : 14] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[258:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[220:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8}}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[205:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8}}}};
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[14 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[220 : 15] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[205:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[200:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8}}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_sums_0[194:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[191 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8}}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 6);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[5 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[200 : 6] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[194:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 20);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[19 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[220 : 20] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[200:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 52);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[51 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[272 : 52] = adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[220:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[127 : 64];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[189 : 128];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19},{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[182:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 7);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[6 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[189 : 7] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[182:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[166:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = NAFElements_sums_0[150:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 16);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[15 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[166 : 16] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[150:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 23);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[22 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[189 : 23] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[166:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[145:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[141:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9}}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 4);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[145 : 4] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[141:0];
  end

  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[129:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[127 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19,{{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9}}};
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[125:0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[125 : 64];
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16},{_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9}};
  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 4);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[3 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[129 : 4] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[125:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 16);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[15 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[145 : 16] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[129:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 44);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p[43 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p[189 : 44] = adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[145:0];
  end

  assign adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 83);
  always @(*) begin
    adder_negMUL_multiElements_lsbMUL_p[82 : 0] = _zz_adder_negMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_lsbMUL_p[272 : 83] = adder_negMUL_multiElements_lsbMUL_multiElements_add_add_io_s[189:0];
  end

  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = NAFElements_sums_0[120:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[96:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10}};
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[23 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[120 : 24] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[96:0];
  end

  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[84:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[74:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10}};
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 10);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[9 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[84 : 10] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[74:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 36);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[35 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[120 : 36] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[84:0];
  end

  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[68:0];
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14,{_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10}};
  assign _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 0];
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p = {_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5,_zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9};
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 5);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[68 : 5] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[63:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 4);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[3 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[58 : 4] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[54:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 10);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[9 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[68 : 10] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_add_add_io_s[58:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 52);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p[51 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p[120 : 52] = adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_add_add_io_s[68:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p = _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
  assign adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p = _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p[26 : 0] = _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p[36 : 27] = adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_add_add_io_s[9:0];
  end

  assign adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 84);
  always @(*) begin
    adder_negMUL_multiElements_msbMUL_p[83 : 0] = _zz_adder_negMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_p[120 : 84] = adder_negMUL_multiElements_msbMUL_multiElements_add_add_io_s[36:0];
  end

  assign adder_negMUL_multiElements_add_add_io_a = (adder_negMUL_multiElements_lsbMUL_p >>> 152);
  always @(*) begin
    adder_negMUL_p[151 : 0] = _zz_adder_negMUL_p;
    adder_negMUL_p[272 : 152] = adder_negMUL_multiElements_add_add_io_s[120:0];
  end

  assign adder_add_io_b = ({106'd0,adder_negMUL_p_delay_1} <<< 106);
  assign io_p[378 : 0] = _zz_io_p;
  always @(posedge clk) begin
    _zz_NAFElements_sums_0_1 <= _zz_NAFElements_sums_0[127 : 64];
    _zz_NAFElements_sums_0_2 <= _zz_NAFElements_sums_0[191 : 128];
    _zz_NAFElements_sums_0_3 <= _zz_NAFElements_sums_0_2;
    _zz_NAFElements_sums_0_4 <= _zz_NAFElements_sums_0[255 : 192];
    _zz_NAFElements_sums_0_5 <= _zz_NAFElements_sums_0_4;
    _zz_NAFElements_sums_0_6 <= _zz_NAFElements_sums_0_5;
    _zz_NAFElements_sums_0_7 <= _zz_NAFElements_sums_0[319 : 256];
    _zz_NAFElements_sums_0_8 <= _zz_NAFElements_sums_0_7;
    _zz_NAFElements_sums_0_9 <= _zz_NAFElements_sums_0_8;
    _zz_NAFElements_sums_0_10 <= _zz_NAFElements_sums_0_9;
    _zz_NAFElements_sums_0_11 <= _zz_NAFElements_sums_0[378 : 320];
    _zz_NAFElements_sums_0_12 <= _zz_NAFElements_sums_0_11;
    _zz_NAFElements_sums_0_13 <= _zz_NAFElements_sums_0_12;
    _zz_NAFElements_sums_0_14 <= _zz_NAFElements_sums_0_13;
    _zz_NAFElements_sums_0_15 <= _zz_NAFElements_sums_0_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 18];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 18];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[63 : 18];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5[63 : 18];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6[63 : 18];
    _zz_io_a <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 46);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[45 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5[63 : 13];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 8];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 8];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4[63 : 8];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5[63 : 8];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6[63 : 8];
    _zz_io_a_1 <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 5);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[50 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[63 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5[59 : 1];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 36];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[35 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 36];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[35 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 36];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[35 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[63 : 36];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[35 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[286 : 256];
    _zz_io_a_2 <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 29);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[28 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 30];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[29 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 30];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[29 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 30];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[29 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[63 : 30];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[29 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[280 : 256];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 26];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 26];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 26];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4[63 : 26];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[276 : 256];
    _zz_io_a_3 <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 4);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[34 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[62 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 12];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[11 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 12];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[11 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 12];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[11 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[63 : 12];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[11 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[262 : 256];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 3];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[2 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 3];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[2 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 3];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[2 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[61 : 3];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[2 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[8 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 53];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[52 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 53];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[52 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 53];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[52 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[239 : 192];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[234 : 192];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_io_a_4 <= (adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 23);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[22 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 28];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[27 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 28];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[27 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 28];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[27 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[214 : 192];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 23];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[22 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 23];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[22 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 23];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[22 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[209 : 192];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
    adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1 <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 54];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[53 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 54];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[53 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[176 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[170 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[5 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[37 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[115 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 40];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[39 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 40];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[39 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[162 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 32];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[31 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 32];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[31 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[154 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
    _zz_io_a_5 <= (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 8);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[7 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 14];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[13 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 14];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[13 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[136 : 128];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 58];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[57 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[116 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[19 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 53];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[52 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[111 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 48];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[106 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1 <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 43];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[42 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[101 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 33];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[32 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[91 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
    adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1 <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[9 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[9 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[50 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 21];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[20 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[79 : 64];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[50 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[28 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[46 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[42 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_io_a_6 <= (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 4);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_io_a_7 <= (adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 33);
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[32 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[31 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[25 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[5 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[20 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[15 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[10 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[47 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[82 : 0];
    _zz_adder_posMUL_multiElements_lsbMUL_p <= adder_posMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[215 : 0];
    _zz_adder_posMUL_multiElements_msbMUL_p <= _zz__zz_adder_posMUL_multiElements_msbMUL_p[4 : 0];
    _zz_adder_posMUL_multiElements_msbMUL_p_1 <= _zz_adder_posMUL_multiElements_msbMUL_p;
    _zz_adder_posMUL_multiElements_msbMUL_p_2 <= _zz_adder_posMUL_multiElements_msbMUL_p_1;
    _zz_adder_posMUL_multiElements_msbMUL_p_3 <= _zz_adder_posMUL_multiElements_msbMUL_p_2;
    _zz_adder_posMUL_multiElements_msbMUL_p_4 <= _zz_adder_posMUL_multiElements_msbMUL_p_3;
    adder_posMUL_multiElements_msbMUL_p_delay_1 <= adder_posMUL_multiElements_msbMUL_p;
    adder_posMUL_multiElements_msbMUL_p_delay_2 <= adder_posMUL_multiElements_msbMUL_p_delay_1;
    adder_posMUL_multiElements_msbMUL_p_delay_3 <= adder_posMUL_multiElements_msbMUL_p_delay_2;
    adder_posMUL_multiElements_msbMUL_p_delay_4 <= adder_posMUL_multiElements_msbMUL_p_delay_3;
    adder_posMUL_multiElements_msbMUL_p_delay_5 <= adder_posMUL_multiElements_msbMUL_p_delay_4;
    _zz_adder_posMUL_p <= adder_posMUL_multiElements_lsbMUL_p[373 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 22];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[21 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 22];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[21 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[63 : 22];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[21 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5[63 : 22];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5[21 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[272 : 256];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 17];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[16 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 17];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[16 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 17];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[16 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[63 : 17];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4[16 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[267 : 256];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[258 : 256];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 39];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[38 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 39];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[38 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 39];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[38 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[225 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[32 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[13 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 34];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[33 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 34];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[33 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 34];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[33 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[220 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[205 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19;
    _zz_io_a_8 <= (adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 15);
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[14 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 14];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[13 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 14];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[13 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[63 : 14];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3[13 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[200 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[63 : 8];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3[7 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[194 : 192];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_20 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19;
    adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1 <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[5 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[19 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[51 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[63 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[61 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 60];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[59 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 60];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[59 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[182 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[6 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 44];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[43 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 44];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[43 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[166 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 28];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[27 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[63 : 28];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[27 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[150 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[15 : 0];
    adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_delay_1 <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[22 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 23];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[22 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[63 : 23];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2[22 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[145 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[63 : 19];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2[18 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[141 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 7];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[6 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[63 : 7];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2[6 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[129 : 128];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_17;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_19 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_18;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[61 : 3];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2[2 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_16 <= _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_15;
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[15 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[43 : 0];
    _zz_adder_negMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[82 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 62];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[61 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[120 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[63 : 38];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1[37 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[96 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_13;
    _zz_io_a_9 <= (adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p >>> 24);
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[23 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[63 : 26];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1[25 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[84 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[63 : 16];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1[15 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p[74 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p_13;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[9 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[35 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[63 : 10];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_5;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_1[9 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_10 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_9;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[68 : 64];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_11;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_12;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_14 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p_13;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[63 : 5];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_5 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_4;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p[4 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_6;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_7;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_9 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p_8;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[4 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[58 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[54 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1 <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[3 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[9 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_multiElements_lsbMUL_p[51 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p <= _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[36 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p_3;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p <= _zz__zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p[9 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_1;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_2;
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_4 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_msbMUL_p_3;
    _zz_io_a_10 <= (adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p >>> 27);
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_multiElements_lsbMUL_p[26 : 0];
    _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_1 <= _zz_adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1 <= adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p;
    adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_2 <= adder_negMUL_multiElements_msbMUL_multiElements_msbMUL_p_delay_1;
    _zz_adder_negMUL_multiElements_msbMUL_p <= adder_negMUL_multiElements_msbMUL_multiElements_lsbMUL_p[83 : 0];
    _zz_adder_negMUL_p <= adder_negMUL_multiElements_lsbMUL_p[151 : 0];
    adder_negMUL_p_delay_1 <= adder_negMUL_p;
  end


endmodule

module KaratsubaMUL_17 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  output     [755:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [47:0]   core_io_a_0;
  wire       [47:0]   core_io_a_1;
  wire       [47:0]   core_io_a_2;
  wire       [47:0]   core_io_a_3;
  wire       [47:0]   core_io_a_4;
  wire       [47:0]   core_io_a_5;
  wire       [47:0]   core_io_a_6;
  wire       [47:0]   core_io_a_7;
  wire       [47:0]   core_io_b_0;
  wire       [47:0]   core_io_b_1;
  wire       [47:0]   core_io_b_2;
  wire       [47:0]   core_io_b_3;
  wire       [47:0]   core_io_b_4;
  wire       [47:0]   core_io_b_5;
  wire       [47:0]   core_io_b_6;
  wire       [47:0]   core_io_b_7;
  wire       [767:0]  core_io_p;
  wire       [47:0]   _zz_io_p_121;
  wire       [239:0]  _zz_io_p_122;
  wire       [383:0]  a;
  wire       [383:0]  b;
  wire       [335:0]  _zz_io_a_0;
  wire       [335:0]  _zz_io_b_0;
  wire       [755:0]  _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;
  reg        [47:0]   _zz_io_p_4;
  reg        [47:0]   _zz_io_p_5;
  reg        [47:0]   _zz_io_p_6;
  reg        [47:0]   _zz_io_p_7;
  reg        [47:0]   _zz_io_p_8;
  reg        [47:0]   _zz_io_p_9;
  reg        [47:0]   _zz_io_p_10;
  reg        [47:0]   _zz_io_p_11;
  reg        [47:0]   _zz_io_p_12;
  reg        [47:0]   _zz_io_p_13;
  reg        [47:0]   _zz_io_p_14;
  reg        [47:0]   _zz_io_p_15;
  reg        [47:0]   _zz_io_p_16;
  reg        [47:0]   _zz_io_p_17;
  reg        [47:0]   _zz_io_p_18;
  reg        [47:0]   _zz_io_p_19;
  reg        [47:0]   _zz_io_p_20;
  reg        [47:0]   _zz_io_p_21;
  reg        [47:0]   _zz_io_p_22;
  reg        [47:0]   _zz_io_p_23;
  reg        [47:0]   _zz_io_p_24;
  reg        [47:0]   _zz_io_p_25;
  reg        [47:0]   _zz_io_p_26;
  reg        [47:0]   _zz_io_p_27;
  reg        [47:0]   _zz_io_p_28;
  reg        [47:0]   _zz_io_p_29;
  reg        [47:0]   _zz_io_p_30;
  reg        [47:0]   _zz_io_p_31;
  reg        [47:0]   _zz_io_p_32;
  reg        [47:0]   _zz_io_p_33;
  reg        [47:0]   _zz_io_p_34;
  reg        [47:0]   _zz_io_p_35;
  reg        [47:0]   _zz_io_p_36;
  reg        [47:0]   _zz_io_p_37;
  reg        [47:0]   _zz_io_p_38;
  reg        [47:0]   _zz_io_p_39;
  reg        [47:0]   _zz_io_p_40;
  reg        [47:0]   _zz_io_p_41;
  reg        [47:0]   _zz_io_p_42;
  reg        [47:0]   _zz_io_p_43;
  reg        [47:0]   _zz_io_p_44;
  reg        [47:0]   _zz_io_p_45;
  reg        [47:0]   _zz_io_p_46;
  reg        [47:0]   _zz_io_p_47;
  reg        [47:0]   _zz_io_p_48;
  reg        [47:0]   _zz_io_p_49;
  reg        [47:0]   _zz_io_p_50;
  reg        [47:0]   _zz_io_p_51;
  reg        [47:0]   _zz_io_p_52;
  reg        [47:0]   _zz_io_p_53;
  reg        [47:0]   _zz_io_p_54;
  reg        [47:0]   _zz_io_p_55;
  reg        [47:0]   _zz_io_p_56;
  reg        [47:0]   _zz_io_p_57;
  reg        [47:0]   _zz_io_p_58;
  reg        [47:0]   _zz_io_p_59;
  reg        [47:0]   _zz_io_p_60;
  reg        [47:0]   _zz_io_p_61;
  reg        [47:0]   _zz_io_p_62;
  reg        [47:0]   _zz_io_p_63;
  reg        [47:0]   _zz_io_p_64;
  reg        [47:0]   _zz_io_p_65;
  reg        [47:0]   _zz_io_p_66;
  reg        [47:0]   _zz_io_p_67;
  reg        [47:0]   _zz_io_p_68;
  reg        [47:0]   _zz_io_p_69;
  reg        [47:0]   _zz_io_p_70;
  reg        [47:0]   _zz_io_p_71;
  reg        [47:0]   _zz_io_p_72;
  reg        [47:0]   _zz_io_p_73;
  reg        [47:0]   _zz_io_p_74;
  reg        [47:0]   _zz_io_p_75;
  reg        [47:0]   _zz_io_p_76;
  reg        [47:0]   _zz_io_p_77;
  reg        [47:0]   _zz_io_p_78;
  reg        [47:0]   _zz_io_p_79;
  reg        [47:0]   _zz_io_p_80;
  reg        [47:0]   _zz_io_p_81;
  reg        [47:0]   _zz_io_p_82;
  reg        [47:0]   _zz_io_p_83;
  reg        [47:0]   _zz_io_p_84;
  reg        [47:0]   _zz_io_p_85;
  reg        [47:0]   _zz_io_p_86;
  reg        [47:0]   _zz_io_p_87;
  reg        [47:0]   _zz_io_p_88;
  reg        [47:0]   _zz_io_p_89;
  reg        [47:0]   _zz_io_p_90;
  reg        [47:0]   _zz_io_p_91;
  reg        [47:0]   _zz_io_p_92;
  reg        [47:0]   _zz_io_p_93;
  reg        [47:0]   _zz_io_p_94;
  reg        [47:0]   _zz_io_p_95;
  reg        [47:0]   _zz_io_p_96;
  reg        [47:0]   _zz_io_p_97;
  reg        [47:0]   _zz_io_p_98;
  reg        [47:0]   _zz_io_p_99;
  reg        [47:0]   _zz_io_p_100;
  reg        [47:0]   _zz_io_p_101;
  reg        [47:0]   _zz_io_p_102;
  reg        [47:0]   _zz_io_p_103;
  reg        [47:0]   _zz_io_p_104;
  reg        [47:0]   _zz_io_p_105;
  reg        [47:0]   _zz_io_p_106;
  reg        [47:0]   _zz_io_p_107;
  reg        [47:0]   _zz_io_p_108;
  reg        [47:0]   _zz_io_p_109;
  reg        [47:0]   _zz_io_p_110;
  reg        [47:0]   _zz_io_p_111;
  reg        [47:0]   _zz_io_p_112;
  reg        [47:0]   _zz_io_p_113;
  reg        [47:0]   _zz_io_p_114;
  reg        [47:0]   _zz_io_p_115;
  reg        [47:0]   _zz_io_p_116;
  reg        [47:0]   _zz_io_p_117;
  reg        [47:0]   _zz_io_p_118;
  reg        [47:0]   _zz_io_p_119;
  reg        [47:0]   _zz_io_p_120;

  assign _zz_io_p_121 = _zz_io_p_75;
  assign _zz_io_p_122 = {_zz_io_p_65,{_zz_io_p_54,{_zz_io_p_42,{_zz_io_p_29,_zz_io_p_15}}}};
  KaratsubaCore_17 core (
    .io_a_0 (core_io_a_0[47:0]), //i
    .io_a_1 (core_io_a_1[47:0]), //i
    .io_a_2 (core_io_a_2[47:0]), //i
    .io_a_3 (core_io_a_3[47:0]), //i
    .io_a_4 (core_io_a_4[47:0]), //i
    .io_a_5 (core_io_a_5[47:0]), //i
    .io_a_6 (core_io_a_6[47:0]), //i
    .io_a_7 (core_io_a_7[47:0]), //i
    .io_b_0 (core_io_b_0[47:0]), //i
    .io_b_1 (core_io_b_1[47:0]), //i
    .io_b_2 (core_io_b_2[47:0]), //i
    .io_b_3 (core_io_b_3[47:0]), //i
    .io_b_4 (core_io_b_4[47:0]), //i
    .io_b_5 (core_io_b_5[47:0]), //i
    .io_b_6 (core_io_b_6[47:0]), //i
    .io_b_7 (core_io_b_7[47:0]), //i
    .io_p   (core_io_p[767:0] ), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  assign a = {6'd0, io_a};
  assign b = {6'd0, io_b};
  assign _zz_io_a_0 = a[335:0];
  assign core_io_a_0 = _zz_io_a_0[47 : 0];
  assign core_io_a_1 = _zz_io_a_0[95 : 48];
  assign core_io_a_2 = _zz_io_a_0[143 : 96];
  assign core_io_a_3 = _zz_io_a_0[191 : 144];
  assign core_io_a_4 = _zz_io_a_0[239 : 192];
  assign core_io_a_5 = _zz_io_a_0[287 : 240];
  assign core_io_a_6 = _zz_io_a_0[335 : 288];
  assign core_io_a_7 = (a >>> 336);
  assign _zz_io_b_0 = b[335:0];
  assign core_io_b_0 = _zz_io_b_0[47 : 0];
  assign core_io_b_1 = _zz_io_b_0[95 : 48];
  assign core_io_b_2 = _zz_io_b_0[143 : 96];
  assign core_io_b_3 = _zz_io_b_0[191 : 144];
  assign core_io_b_4 = _zz_io_b_0[239 : 192];
  assign core_io_b_5 = _zz_io_b_0[287 : 240];
  assign core_io_b_6 = _zz_io_b_0[335 : 288];
  assign core_io_b_7 = (b >>> 336);
  assign _zz_io_p = core_io_p[755:0];
  assign io_p = {_zz_io_p[755 : 720],{_zz_io_p_120,{_zz_io_p_119,{_zz_io_p_117,{_zz_io_p_114,{_zz_io_p_110,{_zz_io_p_105,{_zz_io_p_99,{_zz_io_p_92,{_zz_io_p_84,{_zz_io_p_121,_zz_io_p_122}}}}}}}}}}};
  always @(posedge clk) begin
    _zz_io_p_1 <= _zz_io_p[47 : 0];
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= _zz_io_p_2;
    _zz_io_p_4 <= _zz_io_p_3;
    _zz_io_p_5 <= _zz_io_p_4;
    _zz_io_p_6 <= _zz_io_p_5;
    _zz_io_p_7 <= _zz_io_p_6;
    _zz_io_p_8 <= _zz_io_p_7;
    _zz_io_p_9 <= _zz_io_p_8;
    _zz_io_p_10 <= _zz_io_p_9;
    _zz_io_p_11 <= _zz_io_p_10;
    _zz_io_p_12 <= _zz_io_p_11;
    _zz_io_p_13 <= _zz_io_p_12;
    _zz_io_p_14 <= _zz_io_p_13;
    _zz_io_p_15 <= _zz_io_p_14;
    _zz_io_p_16 <= _zz_io_p[95 : 48];
    _zz_io_p_17 <= _zz_io_p_16;
    _zz_io_p_18 <= _zz_io_p_17;
    _zz_io_p_19 <= _zz_io_p_18;
    _zz_io_p_20 <= _zz_io_p_19;
    _zz_io_p_21 <= _zz_io_p_20;
    _zz_io_p_22 <= _zz_io_p_21;
    _zz_io_p_23 <= _zz_io_p_22;
    _zz_io_p_24 <= _zz_io_p_23;
    _zz_io_p_25 <= _zz_io_p_24;
    _zz_io_p_26 <= _zz_io_p_25;
    _zz_io_p_27 <= _zz_io_p_26;
    _zz_io_p_28 <= _zz_io_p_27;
    _zz_io_p_29 <= _zz_io_p_28;
    _zz_io_p_30 <= _zz_io_p[143 : 96];
    _zz_io_p_31 <= _zz_io_p_30;
    _zz_io_p_32 <= _zz_io_p_31;
    _zz_io_p_33 <= _zz_io_p_32;
    _zz_io_p_34 <= _zz_io_p_33;
    _zz_io_p_35 <= _zz_io_p_34;
    _zz_io_p_36 <= _zz_io_p_35;
    _zz_io_p_37 <= _zz_io_p_36;
    _zz_io_p_38 <= _zz_io_p_37;
    _zz_io_p_39 <= _zz_io_p_38;
    _zz_io_p_40 <= _zz_io_p_39;
    _zz_io_p_41 <= _zz_io_p_40;
    _zz_io_p_42 <= _zz_io_p_41;
    _zz_io_p_43 <= _zz_io_p[191 : 144];
    _zz_io_p_44 <= _zz_io_p_43;
    _zz_io_p_45 <= _zz_io_p_44;
    _zz_io_p_46 <= _zz_io_p_45;
    _zz_io_p_47 <= _zz_io_p_46;
    _zz_io_p_48 <= _zz_io_p_47;
    _zz_io_p_49 <= _zz_io_p_48;
    _zz_io_p_50 <= _zz_io_p_49;
    _zz_io_p_51 <= _zz_io_p_50;
    _zz_io_p_52 <= _zz_io_p_51;
    _zz_io_p_53 <= _zz_io_p_52;
    _zz_io_p_54 <= _zz_io_p_53;
    _zz_io_p_55 <= _zz_io_p[239 : 192];
    _zz_io_p_56 <= _zz_io_p_55;
    _zz_io_p_57 <= _zz_io_p_56;
    _zz_io_p_58 <= _zz_io_p_57;
    _zz_io_p_59 <= _zz_io_p_58;
    _zz_io_p_60 <= _zz_io_p_59;
    _zz_io_p_61 <= _zz_io_p_60;
    _zz_io_p_62 <= _zz_io_p_61;
    _zz_io_p_63 <= _zz_io_p_62;
    _zz_io_p_64 <= _zz_io_p_63;
    _zz_io_p_65 <= _zz_io_p_64;
    _zz_io_p_66 <= _zz_io_p[287 : 240];
    _zz_io_p_67 <= _zz_io_p_66;
    _zz_io_p_68 <= _zz_io_p_67;
    _zz_io_p_69 <= _zz_io_p_68;
    _zz_io_p_70 <= _zz_io_p_69;
    _zz_io_p_71 <= _zz_io_p_70;
    _zz_io_p_72 <= _zz_io_p_71;
    _zz_io_p_73 <= _zz_io_p_72;
    _zz_io_p_74 <= _zz_io_p_73;
    _zz_io_p_75 <= _zz_io_p_74;
    _zz_io_p_76 <= _zz_io_p[335 : 288];
    _zz_io_p_77 <= _zz_io_p_76;
    _zz_io_p_78 <= _zz_io_p_77;
    _zz_io_p_79 <= _zz_io_p_78;
    _zz_io_p_80 <= _zz_io_p_79;
    _zz_io_p_81 <= _zz_io_p_80;
    _zz_io_p_82 <= _zz_io_p_81;
    _zz_io_p_83 <= _zz_io_p_82;
    _zz_io_p_84 <= _zz_io_p_83;
    _zz_io_p_85 <= _zz_io_p[383 : 336];
    _zz_io_p_86 <= _zz_io_p_85;
    _zz_io_p_87 <= _zz_io_p_86;
    _zz_io_p_88 <= _zz_io_p_87;
    _zz_io_p_89 <= _zz_io_p_88;
    _zz_io_p_90 <= _zz_io_p_89;
    _zz_io_p_91 <= _zz_io_p_90;
    _zz_io_p_92 <= _zz_io_p_91;
    _zz_io_p_93 <= _zz_io_p[431 : 384];
    _zz_io_p_94 <= _zz_io_p_93;
    _zz_io_p_95 <= _zz_io_p_94;
    _zz_io_p_96 <= _zz_io_p_95;
    _zz_io_p_97 <= _zz_io_p_96;
    _zz_io_p_98 <= _zz_io_p_97;
    _zz_io_p_99 <= _zz_io_p_98;
    _zz_io_p_100 <= _zz_io_p[479 : 432];
    _zz_io_p_101 <= _zz_io_p_100;
    _zz_io_p_102 <= _zz_io_p_101;
    _zz_io_p_103 <= _zz_io_p_102;
    _zz_io_p_104 <= _zz_io_p_103;
    _zz_io_p_105 <= _zz_io_p_104;
    _zz_io_p_106 <= _zz_io_p[527 : 480];
    _zz_io_p_107 <= _zz_io_p_106;
    _zz_io_p_108 <= _zz_io_p_107;
    _zz_io_p_109 <= _zz_io_p_108;
    _zz_io_p_110 <= _zz_io_p_109;
    _zz_io_p_111 <= _zz_io_p[575 : 528];
    _zz_io_p_112 <= _zz_io_p_111;
    _zz_io_p_113 <= _zz_io_p_112;
    _zz_io_p_114 <= _zz_io_p_113;
    _zz_io_p_115 <= _zz_io_p[623 : 576];
    _zz_io_p_116 <= _zz_io_p_115;
    _zz_io_p_117 <= _zz_io_p_116;
    _zz_io_p_118 <= _zz_io_p[671 : 624];
    _zz_io_p_119 <= _zz_io_p_118;
    _zz_io_p_120 <= _zz_io_p[719 : 672];
  end


endmodule

module KaratsubaMUL_16 (
  input      [376:0]  io_a,
  input      [376:0]  io_b,
  output     [753:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [47:0]   core_io_a_0;
  wire       [47:0]   core_io_a_1;
  wire       [47:0]   core_io_a_2;
  wire       [47:0]   core_io_a_3;
  wire       [47:0]   core_io_a_4;
  wire       [47:0]   core_io_a_5;
  wire       [47:0]   core_io_a_6;
  wire       [47:0]   core_io_a_7;
  wire       [47:0]   core_io_b_0;
  wire       [47:0]   core_io_b_1;
  wire       [47:0]   core_io_b_2;
  wire       [47:0]   core_io_b_3;
  wire       [47:0]   core_io_b_4;
  wire       [47:0]   core_io_b_5;
  wire       [47:0]   core_io_b_6;
  wire       [47:0]   core_io_b_7;
  wire       [767:0]  core_io_p;
  wire       [47:0]   _zz_io_p_121;
  wire       [239:0]  _zz_io_p_122;
  wire       [383:0]  a;
  wire       [383:0]  b;
  wire       [335:0]  _zz_io_a_0;
  wire       [335:0]  _zz_io_b_0;
  wire       [753:0]  _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;
  reg        [47:0]   _zz_io_p_4;
  reg        [47:0]   _zz_io_p_5;
  reg        [47:0]   _zz_io_p_6;
  reg        [47:0]   _zz_io_p_7;
  reg        [47:0]   _zz_io_p_8;
  reg        [47:0]   _zz_io_p_9;
  reg        [47:0]   _zz_io_p_10;
  reg        [47:0]   _zz_io_p_11;
  reg        [47:0]   _zz_io_p_12;
  reg        [47:0]   _zz_io_p_13;
  reg        [47:0]   _zz_io_p_14;
  reg        [47:0]   _zz_io_p_15;
  reg        [47:0]   _zz_io_p_16;
  reg        [47:0]   _zz_io_p_17;
  reg        [47:0]   _zz_io_p_18;
  reg        [47:0]   _zz_io_p_19;
  reg        [47:0]   _zz_io_p_20;
  reg        [47:0]   _zz_io_p_21;
  reg        [47:0]   _zz_io_p_22;
  reg        [47:0]   _zz_io_p_23;
  reg        [47:0]   _zz_io_p_24;
  reg        [47:0]   _zz_io_p_25;
  reg        [47:0]   _zz_io_p_26;
  reg        [47:0]   _zz_io_p_27;
  reg        [47:0]   _zz_io_p_28;
  reg        [47:0]   _zz_io_p_29;
  reg        [47:0]   _zz_io_p_30;
  reg        [47:0]   _zz_io_p_31;
  reg        [47:0]   _zz_io_p_32;
  reg        [47:0]   _zz_io_p_33;
  reg        [47:0]   _zz_io_p_34;
  reg        [47:0]   _zz_io_p_35;
  reg        [47:0]   _zz_io_p_36;
  reg        [47:0]   _zz_io_p_37;
  reg        [47:0]   _zz_io_p_38;
  reg        [47:0]   _zz_io_p_39;
  reg        [47:0]   _zz_io_p_40;
  reg        [47:0]   _zz_io_p_41;
  reg        [47:0]   _zz_io_p_42;
  reg        [47:0]   _zz_io_p_43;
  reg        [47:0]   _zz_io_p_44;
  reg        [47:0]   _zz_io_p_45;
  reg        [47:0]   _zz_io_p_46;
  reg        [47:0]   _zz_io_p_47;
  reg        [47:0]   _zz_io_p_48;
  reg        [47:0]   _zz_io_p_49;
  reg        [47:0]   _zz_io_p_50;
  reg        [47:0]   _zz_io_p_51;
  reg        [47:0]   _zz_io_p_52;
  reg        [47:0]   _zz_io_p_53;
  reg        [47:0]   _zz_io_p_54;
  reg        [47:0]   _zz_io_p_55;
  reg        [47:0]   _zz_io_p_56;
  reg        [47:0]   _zz_io_p_57;
  reg        [47:0]   _zz_io_p_58;
  reg        [47:0]   _zz_io_p_59;
  reg        [47:0]   _zz_io_p_60;
  reg        [47:0]   _zz_io_p_61;
  reg        [47:0]   _zz_io_p_62;
  reg        [47:0]   _zz_io_p_63;
  reg        [47:0]   _zz_io_p_64;
  reg        [47:0]   _zz_io_p_65;
  reg        [47:0]   _zz_io_p_66;
  reg        [47:0]   _zz_io_p_67;
  reg        [47:0]   _zz_io_p_68;
  reg        [47:0]   _zz_io_p_69;
  reg        [47:0]   _zz_io_p_70;
  reg        [47:0]   _zz_io_p_71;
  reg        [47:0]   _zz_io_p_72;
  reg        [47:0]   _zz_io_p_73;
  reg        [47:0]   _zz_io_p_74;
  reg        [47:0]   _zz_io_p_75;
  reg        [47:0]   _zz_io_p_76;
  reg        [47:0]   _zz_io_p_77;
  reg        [47:0]   _zz_io_p_78;
  reg        [47:0]   _zz_io_p_79;
  reg        [47:0]   _zz_io_p_80;
  reg        [47:0]   _zz_io_p_81;
  reg        [47:0]   _zz_io_p_82;
  reg        [47:0]   _zz_io_p_83;
  reg        [47:0]   _zz_io_p_84;
  reg        [47:0]   _zz_io_p_85;
  reg        [47:0]   _zz_io_p_86;
  reg        [47:0]   _zz_io_p_87;
  reg        [47:0]   _zz_io_p_88;
  reg        [47:0]   _zz_io_p_89;
  reg        [47:0]   _zz_io_p_90;
  reg        [47:0]   _zz_io_p_91;
  reg        [47:0]   _zz_io_p_92;
  reg        [47:0]   _zz_io_p_93;
  reg        [47:0]   _zz_io_p_94;
  reg        [47:0]   _zz_io_p_95;
  reg        [47:0]   _zz_io_p_96;
  reg        [47:0]   _zz_io_p_97;
  reg        [47:0]   _zz_io_p_98;
  reg        [47:0]   _zz_io_p_99;
  reg        [47:0]   _zz_io_p_100;
  reg        [47:0]   _zz_io_p_101;
  reg        [47:0]   _zz_io_p_102;
  reg        [47:0]   _zz_io_p_103;
  reg        [47:0]   _zz_io_p_104;
  reg        [47:0]   _zz_io_p_105;
  reg        [47:0]   _zz_io_p_106;
  reg        [47:0]   _zz_io_p_107;
  reg        [47:0]   _zz_io_p_108;
  reg        [47:0]   _zz_io_p_109;
  reg        [47:0]   _zz_io_p_110;
  reg        [47:0]   _zz_io_p_111;
  reg        [47:0]   _zz_io_p_112;
  reg        [47:0]   _zz_io_p_113;
  reg        [47:0]   _zz_io_p_114;
  reg        [47:0]   _zz_io_p_115;
  reg        [47:0]   _zz_io_p_116;
  reg        [47:0]   _zz_io_p_117;
  reg        [47:0]   _zz_io_p_118;
  reg        [47:0]   _zz_io_p_119;
  reg        [47:0]   _zz_io_p_120;

  assign _zz_io_p_121 = _zz_io_p_75;
  assign _zz_io_p_122 = {_zz_io_p_65,{_zz_io_p_54,{_zz_io_p_42,{_zz_io_p_29,_zz_io_p_15}}}};
  KaratsubaCore_17 core (
    .io_a_0 (core_io_a_0[47:0]), //i
    .io_a_1 (core_io_a_1[47:0]), //i
    .io_a_2 (core_io_a_2[47:0]), //i
    .io_a_3 (core_io_a_3[47:0]), //i
    .io_a_4 (core_io_a_4[47:0]), //i
    .io_a_5 (core_io_a_5[47:0]), //i
    .io_a_6 (core_io_a_6[47:0]), //i
    .io_a_7 (core_io_a_7[47:0]), //i
    .io_b_0 (core_io_b_0[47:0]), //i
    .io_b_1 (core_io_b_1[47:0]), //i
    .io_b_2 (core_io_b_2[47:0]), //i
    .io_b_3 (core_io_b_3[47:0]), //i
    .io_b_4 (core_io_b_4[47:0]), //i
    .io_b_5 (core_io_b_5[47:0]), //i
    .io_b_6 (core_io_b_6[47:0]), //i
    .io_b_7 (core_io_b_7[47:0]), //i
    .io_p   (core_io_p[767:0] ), //o
    .clk    (clk              ), //i
    .resetn (resetn           )  //i
  );
  assign a = {7'd0, io_a};
  assign b = {7'd0, io_b};
  assign _zz_io_a_0 = a[335:0];
  assign core_io_a_0 = _zz_io_a_0[47 : 0];
  assign core_io_a_1 = _zz_io_a_0[95 : 48];
  assign core_io_a_2 = _zz_io_a_0[143 : 96];
  assign core_io_a_3 = _zz_io_a_0[191 : 144];
  assign core_io_a_4 = _zz_io_a_0[239 : 192];
  assign core_io_a_5 = _zz_io_a_0[287 : 240];
  assign core_io_a_6 = _zz_io_a_0[335 : 288];
  assign core_io_a_7 = (a >>> 336);
  assign _zz_io_b_0 = b[335:0];
  assign core_io_b_0 = _zz_io_b_0[47 : 0];
  assign core_io_b_1 = _zz_io_b_0[95 : 48];
  assign core_io_b_2 = _zz_io_b_0[143 : 96];
  assign core_io_b_3 = _zz_io_b_0[191 : 144];
  assign core_io_b_4 = _zz_io_b_0[239 : 192];
  assign core_io_b_5 = _zz_io_b_0[287 : 240];
  assign core_io_b_6 = _zz_io_b_0[335 : 288];
  assign core_io_b_7 = (b >>> 336);
  assign _zz_io_p = core_io_p[753:0];
  assign io_p = {_zz_io_p[753 : 720],{_zz_io_p_120,{_zz_io_p_119,{_zz_io_p_117,{_zz_io_p_114,{_zz_io_p_110,{_zz_io_p_105,{_zz_io_p_99,{_zz_io_p_92,{_zz_io_p_84,{_zz_io_p_121,_zz_io_p_122}}}}}}}}}}};
  always @(posedge clk) begin
    _zz_io_p_1 <= _zz_io_p[47 : 0];
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= _zz_io_p_2;
    _zz_io_p_4 <= _zz_io_p_3;
    _zz_io_p_5 <= _zz_io_p_4;
    _zz_io_p_6 <= _zz_io_p_5;
    _zz_io_p_7 <= _zz_io_p_6;
    _zz_io_p_8 <= _zz_io_p_7;
    _zz_io_p_9 <= _zz_io_p_8;
    _zz_io_p_10 <= _zz_io_p_9;
    _zz_io_p_11 <= _zz_io_p_10;
    _zz_io_p_12 <= _zz_io_p_11;
    _zz_io_p_13 <= _zz_io_p_12;
    _zz_io_p_14 <= _zz_io_p_13;
    _zz_io_p_15 <= _zz_io_p_14;
    _zz_io_p_16 <= _zz_io_p[95 : 48];
    _zz_io_p_17 <= _zz_io_p_16;
    _zz_io_p_18 <= _zz_io_p_17;
    _zz_io_p_19 <= _zz_io_p_18;
    _zz_io_p_20 <= _zz_io_p_19;
    _zz_io_p_21 <= _zz_io_p_20;
    _zz_io_p_22 <= _zz_io_p_21;
    _zz_io_p_23 <= _zz_io_p_22;
    _zz_io_p_24 <= _zz_io_p_23;
    _zz_io_p_25 <= _zz_io_p_24;
    _zz_io_p_26 <= _zz_io_p_25;
    _zz_io_p_27 <= _zz_io_p_26;
    _zz_io_p_28 <= _zz_io_p_27;
    _zz_io_p_29 <= _zz_io_p_28;
    _zz_io_p_30 <= _zz_io_p[143 : 96];
    _zz_io_p_31 <= _zz_io_p_30;
    _zz_io_p_32 <= _zz_io_p_31;
    _zz_io_p_33 <= _zz_io_p_32;
    _zz_io_p_34 <= _zz_io_p_33;
    _zz_io_p_35 <= _zz_io_p_34;
    _zz_io_p_36 <= _zz_io_p_35;
    _zz_io_p_37 <= _zz_io_p_36;
    _zz_io_p_38 <= _zz_io_p_37;
    _zz_io_p_39 <= _zz_io_p_38;
    _zz_io_p_40 <= _zz_io_p_39;
    _zz_io_p_41 <= _zz_io_p_40;
    _zz_io_p_42 <= _zz_io_p_41;
    _zz_io_p_43 <= _zz_io_p[191 : 144];
    _zz_io_p_44 <= _zz_io_p_43;
    _zz_io_p_45 <= _zz_io_p_44;
    _zz_io_p_46 <= _zz_io_p_45;
    _zz_io_p_47 <= _zz_io_p_46;
    _zz_io_p_48 <= _zz_io_p_47;
    _zz_io_p_49 <= _zz_io_p_48;
    _zz_io_p_50 <= _zz_io_p_49;
    _zz_io_p_51 <= _zz_io_p_50;
    _zz_io_p_52 <= _zz_io_p_51;
    _zz_io_p_53 <= _zz_io_p_52;
    _zz_io_p_54 <= _zz_io_p_53;
    _zz_io_p_55 <= _zz_io_p[239 : 192];
    _zz_io_p_56 <= _zz_io_p_55;
    _zz_io_p_57 <= _zz_io_p_56;
    _zz_io_p_58 <= _zz_io_p_57;
    _zz_io_p_59 <= _zz_io_p_58;
    _zz_io_p_60 <= _zz_io_p_59;
    _zz_io_p_61 <= _zz_io_p_60;
    _zz_io_p_62 <= _zz_io_p_61;
    _zz_io_p_63 <= _zz_io_p_62;
    _zz_io_p_64 <= _zz_io_p_63;
    _zz_io_p_65 <= _zz_io_p_64;
    _zz_io_p_66 <= _zz_io_p[287 : 240];
    _zz_io_p_67 <= _zz_io_p_66;
    _zz_io_p_68 <= _zz_io_p_67;
    _zz_io_p_69 <= _zz_io_p_68;
    _zz_io_p_70 <= _zz_io_p_69;
    _zz_io_p_71 <= _zz_io_p_70;
    _zz_io_p_72 <= _zz_io_p_71;
    _zz_io_p_73 <= _zz_io_p_72;
    _zz_io_p_74 <= _zz_io_p_73;
    _zz_io_p_75 <= _zz_io_p_74;
    _zz_io_p_76 <= _zz_io_p[335 : 288];
    _zz_io_p_77 <= _zz_io_p_76;
    _zz_io_p_78 <= _zz_io_p_77;
    _zz_io_p_79 <= _zz_io_p_78;
    _zz_io_p_80 <= _zz_io_p_79;
    _zz_io_p_81 <= _zz_io_p_80;
    _zz_io_p_82 <= _zz_io_p_81;
    _zz_io_p_83 <= _zz_io_p_82;
    _zz_io_p_84 <= _zz_io_p_83;
    _zz_io_p_85 <= _zz_io_p[383 : 336];
    _zz_io_p_86 <= _zz_io_p_85;
    _zz_io_p_87 <= _zz_io_p_86;
    _zz_io_p_88 <= _zz_io_p_87;
    _zz_io_p_89 <= _zz_io_p_88;
    _zz_io_p_90 <= _zz_io_p_89;
    _zz_io_p_91 <= _zz_io_p_90;
    _zz_io_p_92 <= _zz_io_p_91;
    _zz_io_p_93 <= _zz_io_p[431 : 384];
    _zz_io_p_94 <= _zz_io_p_93;
    _zz_io_p_95 <= _zz_io_p_94;
    _zz_io_p_96 <= _zz_io_p_95;
    _zz_io_p_97 <= _zz_io_p_96;
    _zz_io_p_98 <= _zz_io_p_97;
    _zz_io_p_99 <= _zz_io_p_98;
    _zz_io_p_100 <= _zz_io_p[479 : 432];
    _zz_io_p_101 <= _zz_io_p_100;
    _zz_io_p_102 <= _zz_io_p_101;
    _zz_io_p_103 <= _zz_io_p_102;
    _zz_io_p_104 <= _zz_io_p_103;
    _zz_io_p_105 <= _zz_io_p_104;
    _zz_io_p_106 <= _zz_io_p[527 : 480];
    _zz_io_p_107 <= _zz_io_p_106;
    _zz_io_p_108 <= _zz_io_p_107;
    _zz_io_p_109 <= _zz_io_p_108;
    _zz_io_p_110 <= _zz_io_p_109;
    _zz_io_p_111 <= _zz_io_p[575 : 528];
    _zz_io_p_112 <= _zz_io_p_111;
    _zz_io_p_113 <= _zz_io_p_112;
    _zz_io_p_114 <= _zz_io_p_113;
    _zz_io_p_115 <= _zz_io_p[623 : 576];
    _zz_io_p_116 <= _zz_io_p_115;
    _zz_io_p_117 <= _zz_io_p_116;
    _zz_io_p_118 <= _zz_io_p[671 : 624];
    _zz_io_p_119 <= _zz_io_p_118;
    _zz_io_p_120 <= _zz_io_p[719 : 672];
  end


endmodule

//BADD_19 replaced by BADD_650

//BADD_20 replaced by BADD_650

//BADD_21 replaced by BADD_650

//BADD_22 replaced by BADD_650

//BADD_23 replaced by BADD_26

//BADD_24 replaced by BADD_26

//BADD_25 replaced by BADD_26

module BADD_26 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  input               io_c,
  output reg [378:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [377:0]  _zz__zz_io_s_1;
  wire       [64:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_8;
  wire       [377:0]  _zz__zz_io_s_8_1;
  wire       [64:0]   _zz__zz_io_s_8_2;
  wire       [0:0]    _zz__zz_io_s_8_3;
  wire       [64:0]   _zz__zz_io_s_15;
  wire       [377:0]  _zz__zz_io_s_15_1;
  wire       [64:0]   _zz__zz_io_s_15_2;
  wire       [0:0]    _zz__zz_io_s_15_3;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [377:0]  _zz__zz_io_s_21_1;
  wire       [64:0]   _zz__zz_io_s_21_2;
  wire       [0:0]    _zz__zz_io_s_21_3;
  wire       [64:0]   _zz__zz_io_s_26;
  wire       [377:0]  _zz__zz_io_s_26_1;
  wire       [64:0]   _zz__zz_io_s_26_2;
  wire       [0:0]    _zz__zz_io_s_26_3;
  wire       [58:0]   _zz__zz_io_s_30;
  wire       [377:0]  _zz__zz_io_s_30_1;
  wire       [58:0]   _zz__zz_io_s_30_2;
  wire       [0:0]    _zz__zz_io_s_30_3;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  wire       [64:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [64:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg                 _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg        [63:0]   _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg                 _zz_io_s_25;
  wire       [64:0]   _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg                 _zz_io_s_29;
  wire       [58:0]   _zz_io_s_30;
  reg        [57:0]   _zz_io_s_31;
  reg                 _zz_io_s_32;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,_zz__zz_io_s_1[63 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {64'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_8 = ({1'b0,io_a[127 : 64]} + {1'b0,_zz__zz_io_s_8_1[127 : 64]});
  assign _zz__zz_io_s_8_1 = (~ io_b);
  assign _zz__zz_io_s_8_3 = _zz_io_s_7;
  assign _zz__zz_io_s_8_2 = {64'd0, _zz__zz_io_s_8_3};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[191 : 128]} + {1'b0,_zz__zz_io_s_15_1[191 : 128]});
  assign _zz__zz_io_s_15_1 = (~ io_b);
  assign _zz__zz_io_s_15_3 = _zz_io_s_14;
  assign _zz__zz_io_s_15_2 = {64'd0, _zz__zz_io_s_15_3};
  assign _zz__zz_io_s_21 = ({1'b0,io_a[255 : 192]} + {1'b0,_zz__zz_io_s_21_1[255 : 192]});
  assign _zz__zz_io_s_21_1 = (~ io_b);
  assign _zz__zz_io_s_21_3 = _zz_io_s_20;
  assign _zz__zz_io_s_21_2 = {64'd0, _zz__zz_io_s_21_3};
  assign _zz__zz_io_s_26 = ({1'b0,io_a[319 : 256]} + {1'b0,_zz__zz_io_s_26_1[319 : 256]});
  assign _zz__zz_io_s_26_1 = (~ io_b);
  assign _zz__zz_io_s_26_3 = _zz_io_s_25;
  assign _zz__zz_io_s_26_2 = {64'd0, _zz__zz_io_s_26_3};
  assign _zz__zz_io_s_30 = ({1'b0,io_a[377 : 320]} + {1'b0,_zz__zz_io_s_30_1[377 : 320]});
  assign _zz__zz_io_s_30_1 = (~ io_b);
  assign _zz__zz_io_s_30_3 = _zz_io_s_29;
  assign _zz__zz_io_s_30_2 = {58'd0, _zz__zz_io_s_30_3};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_6;
    io_s[127 : 64] = _zz_io_s_13;
    io_s[191 : 128] = _zz_io_s_19;
    io_s[255 : 192] = _zz_io_s_24;
    io_s[319 : 256] = _zz_io_s_28;
    io_s[377 : 320] = _zz_io_s_31;
    io_s[378] = (! _zz_io_s_32);
  end

  assign _zz_io_s_8 = (_zz__zz_io_s_8 + _zz__zz_io_s_8_2);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_2);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_2);
  assign _zz_io_s_26 = (_zz__zz_io_s_26 + _zz__zz_io_s_26_2);
  assign _zz_io_s_30 = (_zz__zz_io_s_30 + _zz__zz_io_s_30_2);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= _zz_io_s[64];
    _zz_io_s_9 <= _zz_io_s_8[63:0];
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= _zz_io_s_11;
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_8[64];
    _zz_io_s_16 <= _zz_io_s_15[63:0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_15[64];
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_22;
    _zz_io_s_24 <= _zz_io_s_23;
    _zz_io_s_25 <= _zz_io_s_21[64];
    _zz_io_s_27 <= _zz_io_s_26[63:0];
    _zz_io_s_28 <= _zz_io_s_27;
    _zz_io_s_29 <= _zz_io_s_26[64];
    _zz_io_s_31 <= _zz_io_s_30[57:0];
    _zz_io_s_32 <= _zz_io_s_30[58];
  end


endmodule

//FineReduction_18 replaced by FineReduction_26

//BADD_27 replaced by BADD_531

//BADD_89 replaced by BADD_593

//BADD_88 replaced by BADD_592

//BADD_87 replaced by BADD_591

//BADD_86 replaced by BADD_590

//BADD_85 replaced by BADD_589

//BADD_84 replaced by BADD_588

//BADD_83 replaced by BADD_587

//BADD_82 replaced by BADD_586

//BADD_81 replaced by BADD_585

//BADD_80 replaced by BADD_584

//BADD_79 replaced by BADD_583

//BADD_78 replaced by BADD_582

//BADD_77 replaced by BADD_581

//BADD_76 replaced by BADD_580

//BADD_75 replaced by BADD_579

//BADD_74 replaced by BADD_578

//BADD_73 replaced by BADD_577

//BADD_72 replaced by BADD_576

//BADD_71 replaced by BADD_575

//BADD_70 replaced by BADD_574

//BADD_69 replaced by BADD_573

//BADD_68 replaced by BADD_572

//BADD_67 replaced by BADD_571

//BADD_66 replaced by BADD_570

//BADD_65 replaced by BADD_569

//BADD_64 replaced by BADD_568

//BADD_63 replaced by BADD_567

//BADD_62 replaced by BADD_566

//BADD_61 replaced by BADD_565

//BADD_60 replaced by BADD_564

//BADD_59 replaced by BADD_563

//BADD_58 replaced by BADD_562

//BADD_57 replaced by BADD_561

//BADD_56 replaced by BADD_560

//BADD_55 replaced by BADD_559

//BADD_54 replaced by BADD_558

//BADD_53 replaced by BADD_557

//BADD_52 replaced by BADD_556

//BADD_51 replaced by BADD_555

//BADD_50 replaced by BADD_554

//BADD_49 replaced by BADD_553

//BADD_48 replaced by BADD_552

//BADD_47 replaced by BADD_551

//BADD_46 replaced by BADD_550

//BADD_45 replaced by BADD_549

//BADD_44 replaced by BADD_548

//BADD_43 replaced by BADD_547

//BADD_42 replaced by BADD_546

//BADD_41 replaced by BADD_545

//BADD_40 replaced by BADD_544

//BADD_39 replaced by BADD_543

//BADD_38 replaced by BADD_542

//BADD_37 replaced by BADD_541

//BADD_36 replaced by BADD_540

//BADD_35 replaced by BADD_539

//BADD_34 replaced by BADD_538

//BADD_33 replaced by BADD_537

//BADD_32 replaced by BADD_536

//BADD_31 replaced by BADD_535

//BADD_30 replaced by BADD_534

//BADD_29 replaced by BADD_533

//BADD_28 replaced by BADD_532

//KaratsubaCore replaced by KaratsubaCore_17

//KaratsubaCore_1 replaced by KaratsubaCore_17

//FineReduction_19 replaced by FineReduction_26

//BADD_90 replaced by BADD_531

//BADD_152 replaced by BADD_593

//BADD_151 replaced by BADD_592

//BADD_150 replaced by BADD_591

//BADD_149 replaced by BADD_590

//BADD_148 replaced by BADD_589

//BADD_147 replaced by BADD_588

//BADD_146 replaced by BADD_587

//BADD_145 replaced by BADD_586

//BADD_144 replaced by BADD_585

//BADD_143 replaced by BADD_584

//BADD_142 replaced by BADD_583

//BADD_141 replaced by BADD_582

//BADD_140 replaced by BADD_581

//BADD_139 replaced by BADD_580

//BADD_138 replaced by BADD_579

//BADD_137 replaced by BADD_578

//BADD_136 replaced by BADD_577

//BADD_135 replaced by BADD_576

//BADD_134 replaced by BADD_575

//BADD_133 replaced by BADD_574

//BADD_132 replaced by BADD_573

//BADD_131 replaced by BADD_572

//BADD_130 replaced by BADD_571

//BADD_129 replaced by BADD_570

//BADD_128 replaced by BADD_569

//BADD_127 replaced by BADD_568

//BADD_126 replaced by BADD_567

//BADD_125 replaced by BADD_566

//BADD_124 replaced by BADD_565

//BADD_123 replaced by BADD_564

//BADD_122 replaced by BADD_563

//BADD_121 replaced by BADD_562

//BADD_120 replaced by BADD_561

//BADD_119 replaced by BADD_560

//BADD_118 replaced by BADD_559

//BADD_117 replaced by BADD_558

//BADD_116 replaced by BADD_557

//BADD_115 replaced by BADD_556

//BADD_114 replaced by BADD_555

//BADD_113 replaced by BADD_554

//BADD_112 replaced by BADD_553

//BADD_111 replaced by BADD_552

//BADD_110 replaced by BADD_551

//BADD_109 replaced by BADD_550

//BADD_108 replaced by BADD_549

//BADD_107 replaced by BADD_548

//BADD_106 replaced by BADD_547

//BADD_105 replaced by BADD_546

//BADD_104 replaced by BADD_545

//BADD_103 replaced by BADD_544

//BADD_102 replaced by BADD_543

//BADD_101 replaced by BADD_542

//BADD_100 replaced by BADD_541

//BADD_99 replaced by BADD_540

//BADD_98 replaced by BADD_539

//BADD_97 replaced by BADD_538

//BADD_96 replaced by BADD_537

//BADD_95 replaced by BADD_536

//BADD_94 replaced by BADD_535

//BADD_93 replaced by BADD_534

//BADD_92 replaced by BADD_533

//BADD_91 replaced by BADD_532

//KaratsubaCore_2 replaced by KaratsubaCore_17

//KaratsubaCore_3 replaced by KaratsubaCore_17

//FineReduction_20 replaced by FineReduction_26

//BADD_153 replaced by BADD_531

//BADD_215 replaced by BADD_593

//BADD_214 replaced by BADD_592

//BADD_213 replaced by BADD_591

//BADD_212 replaced by BADD_590

//BADD_211 replaced by BADD_589

//BADD_210 replaced by BADD_588

//BADD_209 replaced by BADD_587

//BADD_208 replaced by BADD_586

//BADD_207 replaced by BADD_585

//BADD_206 replaced by BADD_584

//BADD_205 replaced by BADD_583

//BADD_204 replaced by BADD_582

//BADD_203 replaced by BADD_581

//BADD_202 replaced by BADD_580

//BADD_201 replaced by BADD_579

//BADD_200 replaced by BADD_578

//BADD_199 replaced by BADD_577

//BADD_198 replaced by BADD_576

//BADD_197 replaced by BADD_575

//BADD_196 replaced by BADD_574

//BADD_195 replaced by BADD_573

//BADD_194 replaced by BADD_572

//BADD_193 replaced by BADD_571

//BADD_192 replaced by BADD_570

//BADD_191 replaced by BADD_569

//BADD_190 replaced by BADD_568

//BADD_189 replaced by BADD_567

//BADD_188 replaced by BADD_566

//BADD_187 replaced by BADD_565

//BADD_186 replaced by BADD_564

//BADD_185 replaced by BADD_563

//BADD_184 replaced by BADD_562

//BADD_183 replaced by BADD_561

//BADD_182 replaced by BADD_560

//BADD_181 replaced by BADD_559

//BADD_180 replaced by BADD_558

//BADD_179 replaced by BADD_557

//BADD_178 replaced by BADD_556

//BADD_177 replaced by BADD_555

//BADD_176 replaced by BADD_554

//BADD_175 replaced by BADD_553

//BADD_174 replaced by BADD_552

//BADD_173 replaced by BADD_551

//BADD_172 replaced by BADD_550

//BADD_171 replaced by BADD_549

//BADD_170 replaced by BADD_548

//BADD_169 replaced by BADD_547

//BADD_168 replaced by BADD_546

//BADD_167 replaced by BADD_545

//BADD_166 replaced by BADD_544

//BADD_165 replaced by BADD_543

//BADD_164 replaced by BADD_542

//BADD_163 replaced by BADD_541

//BADD_162 replaced by BADD_540

//BADD_161 replaced by BADD_539

//BADD_160 replaced by BADD_538

//BADD_159 replaced by BADD_537

//BADD_158 replaced by BADD_536

//BADD_157 replaced by BADD_535

//BADD_156 replaced by BADD_534

//BADD_155 replaced by BADD_533

//BADD_154 replaced by BADD_532

//KaratsubaCore_4 replaced by KaratsubaCore_17

//KaratsubaCore_5 replaced by KaratsubaCore_17

//FineReduction_21 replaced by FineReduction_26

//BADD_216 replaced by BADD_531

//BADD_278 replaced by BADD_593

//BADD_277 replaced by BADD_592

//BADD_276 replaced by BADD_591

//BADD_275 replaced by BADD_590

//BADD_274 replaced by BADD_589

//BADD_273 replaced by BADD_588

//BADD_272 replaced by BADD_587

//BADD_271 replaced by BADD_586

//BADD_270 replaced by BADD_585

//BADD_269 replaced by BADD_584

//BADD_268 replaced by BADD_583

//BADD_267 replaced by BADD_582

//BADD_266 replaced by BADD_581

//BADD_265 replaced by BADD_580

//BADD_264 replaced by BADD_579

//BADD_263 replaced by BADD_578

//BADD_262 replaced by BADD_577

//BADD_261 replaced by BADD_576

//BADD_260 replaced by BADD_575

//BADD_259 replaced by BADD_574

//BADD_258 replaced by BADD_573

//BADD_257 replaced by BADD_572

//BADD_256 replaced by BADD_571

//BADD_255 replaced by BADD_570

//BADD_254 replaced by BADD_569

//BADD_253 replaced by BADD_568

//BADD_252 replaced by BADD_567

//BADD_251 replaced by BADD_566

//BADD_250 replaced by BADD_565

//BADD_249 replaced by BADD_564

//BADD_248 replaced by BADD_563

//BADD_247 replaced by BADD_562

//BADD_246 replaced by BADD_561

//BADD_245 replaced by BADD_560

//BADD_244 replaced by BADD_559

//BADD_243 replaced by BADD_558

//BADD_242 replaced by BADD_557

//BADD_241 replaced by BADD_556

//BADD_240 replaced by BADD_555

//BADD_239 replaced by BADD_554

//BADD_238 replaced by BADD_553

//BADD_237 replaced by BADD_552

//BADD_236 replaced by BADD_551

//BADD_235 replaced by BADD_550

//BADD_234 replaced by BADD_549

//BADD_233 replaced by BADD_548

//BADD_232 replaced by BADD_547

//BADD_231 replaced by BADD_546

//BADD_230 replaced by BADD_545

//BADD_229 replaced by BADD_544

//BADD_228 replaced by BADD_543

//BADD_227 replaced by BADD_542

//BADD_226 replaced by BADD_541

//BADD_225 replaced by BADD_540

//BADD_224 replaced by BADD_539

//BADD_223 replaced by BADD_538

//BADD_222 replaced by BADD_537

//BADD_221 replaced by BADD_536

//BADD_220 replaced by BADD_535

//BADD_219 replaced by BADD_534

//BADD_218 replaced by BADD_533

//BADD_217 replaced by BADD_532

//KaratsubaCore_6 replaced by KaratsubaCore_17

//KaratsubaCore_7 replaced by KaratsubaCore_17

//FineReduction_22 replaced by FineReduction_26

//BADD_279 replaced by BADD_531

//BADD_341 replaced by BADD_593

//BADD_340 replaced by BADD_592

//BADD_339 replaced by BADD_591

//BADD_338 replaced by BADD_590

//BADD_337 replaced by BADD_589

//BADD_336 replaced by BADD_588

//BADD_335 replaced by BADD_587

//BADD_334 replaced by BADD_586

//BADD_333 replaced by BADD_585

//BADD_332 replaced by BADD_584

//BADD_331 replaced by BADD_583

//BADD_330 replaced by BADD_582

//BADD_329 replaced by BADD_581

//BADD_328 replaced by BADD_580

//BADD_327 replaced by BADD_579

//BADD_326 replaced by BADD_578

//BADD_325 replaced by BADD_577

//BADD_324 replaced by BADD_576

//BADD_323 replaced by BADD_575

//BADD_322 replaced by BADD_574

//BADD_321 replaced by BADD_573

//BADD_320 replaced by BADD_572

//BADD_319 replaced by BADD_571

//BADD_318 replaced by BADD_570

//BADD_317 replaced by BADD_569

//BADD_316 replaced by BADD_568

//BADD_315 replaced by BADD_567

//BADD_314 replaced by BADD_566

//BADD_313 replaced by BADD_565

//BADD_312 replaced by BADD_564

//BADD_311 replaced by BADD_563

//BADD_310 replaced by BADD_562

//BADD_309 replaced by BADD_561

//BADD_308 replaced by BADD_560

//BADD_307 replaced by BADD_559

//BADD_306 replaced by BADD_558

//BADD_305 replaced by BADD_557

//BADD_304 replaced by BADD_556

//BADD_303 replaced by BADD_555

//BADD_302 replaced by BADD_554

//BADD_301 replaced by BADD_553

//BADD_300 replaced by BADD_552

//BADD_299 replaced by BADD_551

//BADD_298 replaced by BADD_550

//BADD_297 replaced by BADD_549

//BADD_296 replaced by BADD_548

//BADD_295 replaced by BADD_547

//BADD_294 replaced by BADD_546

//BADD_293 replaced by BADD_545

//BADD_292 replaced by BADD_544

//BADD_291 replaced by BADD_543

//BADD_290 replaced by BADD_542

//BADD_289 replaced by BADD_541

//BADD_288 replaced by BADD_540

//BADD_287 replaced by BADD_539

//BADD_286 replaced by BADD_538

//BADD_285 replaced by BADD_537

//BADD_284 replaced by BADD_536

//BADD_283 replaced by BADD_535

//BADD_282 replaced by BADD_534

//BADD_281 replaced by BADD_533

//BADD_280 replaced by BADD_532

//KaratsubaCore_8 replaced by KaratsubaCore_17

//KaratsubaCore_9 replaced by KaratsubaCore_17

//FineReduction_23 replaced by FineReduction_26

//BADD_342 replaced by BADD_531

//BADD_404 replaced by BADD_593

//BADD_403 replaced by BADD_592

//BADD_402 replaced by BADD_591

//BADD_401 replaced by BADD_590

//BADD_400 replaced by BADD_589

//BADD_399 replaced by BADD_588

//BADD_398 replaced by BADD_587

//BADD_397 replaced by BADD_586

//BADD_396 replaced by BADD_585

//BADD_395 replaced by BADD_584

//BADD_394 replaced by BADD_583

//BADD_393 replaced by BADD_582

//BADD_392 replaced by BADD_581

//BADD_391 replaced by BADD_580

//BADD_390 replaced by BADD_579

//BADD_389 replaced by BADD_578

//BADD_388 replaced by BADD_577

//BADD_387 replaced by BADD_576

//BADD_386 replaced by BADD_575

//BADD_385 replaced by BADD_574

//BADD_384 replaced by BADD_573

//BADD_383 replaced by BADD_572

//BADD_382 replaced by BADD_571

//BADD_381 replaced by BADD_570

//BADD_380 replaced by BADD_569

//BADD_379 replaced by BADD_568

//BADD_378 replaced by BADD_567

//BADD_377 replaced by BADD_566

//BADD_376 replaced by BADD_565

//BADD_375 replaced by BADD_564

//BADD_374 replaced by BADD_563

//BADD_373 replaced by BADD_562

//BADD_372 replaced by BADD_561

//BADD_371 replaced by BADD_560

//BADD_370 replaced by BADD_559

//BADD_369 replaced by BADD_558

//BADD_368 replaced by BADD_557

//BADD_367 replaced by BADD_556

//BADD_366 replaced by BADD_555

//BADD_365 replaced by BADD_554

//BADD_364 replaced by BADD_553

//BADD_363 replaced by BADD_552

//BADD_362 replaced by BADD_551

//BADD_361 replaced by BADD_550

//BADD_360 replaced by BADD_549

//BADD_359 replaced by BADD_548

//BADD_358 replaced by BADD_547

//BADD_357 replaced by BADD_546

//BADD_356 replaced by BADD_545

//BADD_355 replaced by BADD_544

//BADD_354 replaced by BADD_543

//BADD_353 replaced by BADD_542

//BADD_352 replaced by BADD_541

//BADD_351 replaced by BADD_540

//BADD_350 replaced by BADD_539

//BADD_349 replaced by BADD_538

//BADD_348 replaced by BADD_537

//BADD_347 replaced by BADD_536

//BADD_346 replaced by BADD_535

//BADD_345 replaced by BADD_534

//BADD_344 replaced by BADD_533

//BADD_343 replaced by BADD_532

//KaratsubaCore_10 replaced by KaratsubaCore_17

//KaratsubaCore_11 replaced by KaratsubaCore_17

//FineReduction_24 replaced by FineReduction_26

//BADD_405 replaced by BADD_531

//BADD_467 replaced by BADD_593

//BADD_466 replaced by BADD_592

//BADD_465 replaced by BADD_591

//BADD_464 replaced by BADD_590

//BADD_463 replaced by BADD_589

//BADD_462 replaced by BADD_588

//BADD_461 replaced by BADD_587

//BADD_460 replaced by BADD_586

//BADD_459 replaced by BADD_585

//BADD_458 replaced by BADD_584

//BADD_457 replaced by BADD_583

//BADD_456 replaced by BADD_582

//BADD_455 replaced by BADD_581

//BADD_454 replaced by BADD_580

//BADD_453 replaced by BADD_579

//BADD_452 replaced by BADD_578

//BADD_451 replaced by BADD_577

//BADD_450 replaced by BADD_576

//BADD_449 replaced by BADD_575

//BADD_448 replaced by BADD_574

//BADD_447 replaced by BADD_573

//BADD_446 replaced by BADD_572

//BADD_445 replaced by BADD_571

//BADD_444 replaced by BADD_570

//BADD_443 replaced by BADD_569

//BADD_442 replaced by BADD_568

//BADD_441 replaced by BADD_567

//BADD_440 replaced by BADD_566

//BADD_439 replaced by BADD_565

//BADD_438 replaced by BADD_564

//BADD_437 replaced by BADD_563

//BADD_436 replaced by BADD_562

//BADD_435 replaced by BADD_561

//BADD_434 replaced by BADD_560

//BADD_433 replaced by BADD_559

//BADD_432 replaced by BADD_558

//BADD_431 replaced by BADD_557

//BADD_430 replaced by BADD_556

//BADD_429 replaced by BADD_555

//BADD_428 replaced by BADD_554

//BADD_427 replaced by BADD_553

//BADD_426 replaced by BADD_552

//BADD_425 replaced by BADD_551

//BADD_424 replaced by BADD_550

//BADD_423 replaced by BADD_549

//BADD_422 replaced by BADD_548

//BADD_421 replaced by BADD_547

//BADD_420 replaced by BADD_546

//BADD_419 replaced by BADD_545

//BADD_418 replaced by BADD_544

//BADD_417 replaced by BADD_543

//BADD_416 replaced by BADD_542

//BADD_415 replaced by BADD_541

//BADD_414 replaced by BADD_540

//BADD_413 replaced by BADD_539

//BADD_412 replaced by BADD_538

//BADD_411 replaced by BADD_537

//BADD_410 replaced by BADD_536

//BADD_409 replaced by BADD_535

//BADD_408 replaced by BADD_534

//BADD_407 replaced by BADD_533

//BADD_406 replaced by BADD_532

//KaratsubaCore_12 replaced by KaratsubaCore_17

//KaratsubaCore_13 replaced by KaratsubaCore_17

//FineReduction_25 replaced by FineReduction_26

//BADD_468 replaced by BADD_531

//BADD_530 replaced by BADD_593

//BADD_529 replaced by BADD_592

//BADD_528 replaced by BADD_591

//BADD_527 replaced by BADD_590

//BADD_526 replaced by BADD_589

//BADD_525 replaced by BADD_588

//BADD_524 replaced by BADD_587

//BADD_523 replaced by BADD_586

//BADD_522 replaced by BADD_585

//BADD_521 replaced by BADD_584

//BADD_520 replaced by BADD_583

//BADD_519 replaced by BADD_582

//BADD_518 replaced by BADD_581

//BADD_517 replaced by BADD_580

//BADD_516 replaced by BADD_579

//BADD_515 replaced by BADD_578

//BADD_514 replaced by BADD_577

//BADD_513 replaced by BADD_576

//BADD_512 replaced by BADD_575

//BADD_511 replaced by BADD_574

//BADD_510 replaced by BADD_573

//BADD_509 replaced by BADD_572

//BADD_508 replaced by BADD_571

//BADD_507 replaced by BADD_570

//BADD_506 replaced by BADD_569

//BADD_505 replaced by BADD_568

//BADD_504 replaced by BADD_567

//BADD_503 replaced by BADD_566

//BADD_502 replaced by BADD_565

//BADD_501 replaced by BADD_564

//BADD_500 replaced by BADD_563

//BADD_499 replaced by BADD_562

//BADD_498 replaced by BADD_561

//BADD_497 replaced by BADD_560

//BADD_496 replaced by BADD_559

//BADD_495 replaced by BADD_558

//BADD_494 replaced by BADD_557

//BADD_493 replaced by BADD_556

//BADD_492 replaced by BADD_555

//BADD_491 replaced by BADD_554

//BADD_490 replaced by BADD_553

//BADD_489 replaced by BADD_552

//BADD_488 replaced by BADD_551

//BADD_487 replaced by BADD_550

//BADD_486 replaced by BADD_549

//BADD_485 replaced by BADD_548

//BADD_484 replaced by BADD_547

//BADD_483 replaced by BADD_546

//BADD_482 replaced by BADD_545

//BADD_481 replaced by BADD_544

//BADD_480 replaced by BADD_543

//BADD_479 replaced by BADD_542

//BADD_478 replaced by BADD_541

//BADD_477 replaced by BADD_540

//BADD_476 replaced by BADD_539

//BADD_475 replaced by BADD_538

//BADD_474 replaced by BADD_537

//BADD_473 replaced by BADD_536

//BADD_472 replaced by BADD_535

//BADD_471 replaced by BADD_534

//BADD_470 replaced by BADD_533

//BADD_469 replaced by BADD_532

//KaratsubaCore_14 replaced by KaratsubaCore_17

//KaratsubaCore_15 replaced by KaratsubaCore_17

module FineReduction_26 (
  input      [377:0]  io_a,
  output     [376:0]  io_r,
  input               clk,
  input               resetn
);

  wire       [378:0]  singleAdd_add_io_s;
  wire       [376:0]  _zz__zz_io_r;
  wire       [376:0]  _zz__zz_io_r_1;
  reg        [63:0]   _zz_singleAdd_a;
  reg        [63:0]   _zz_singleAdd_a_1;
  reg        [63:0]   _zz_singleAdd_a_2;
  reg        [63:0]   _zz_singleAdd_a_3;
  reg        [63:0]   _zz_singleAdd_a_4;
  reg        [63:0]   _zz_singleAdd_a_5;
  reg        [63:0]   _zz_singleAdd_a_6;
  reg        [63:0]   _zz_singleAdd_a_7;
  reg        [63:0]   _zz_singleAdd_a_8;
  reg        [63:0]   _zz_singleAdd_a_9;
  reg        [63:0]   _zz_singleAdd_a_10;
  reg        [63:0]   _zz_singleAdd_a_11;
  reg        [63:0]   _zz_singleAdd_a_12;
  reg        [63:0]   _zz_singleAdd_a_13;
  reg        [63:0]   _zz_singleAdd_a_14;
  reg        [63:0]   _zz_singleAdd_a_15;
  reg        [63:0]   _zz_singleAdd_a_16;
  reg        [63:0]   _zz_singleAdd_a_17;
  reg        [63:0]   _zz_singleAdd_a_18;
  reg        [63:0]   _zz_singleAdd_a_19;
  reg        [57:0]   _zz_singleAdd_a_20;
  wire       [377:0]  singleAdd_a;
  reg        [376:0]  _zz_io_r;

  assign _zz__zz_io_r = singleAdd_add_io_s[376:0];
  assign _zz__zz_io_r_1 = singleAdd_a[376:0];
  BADD_650 singleAdd_add (
    .io_a   (io_a[377:0]                                                                                         ), //i
    .io_b   (378'h1ae3a4617c510eac63b05c06ca1493b1a22d9f300f5138f1ef3622fba094800170b5d44300000008508c00000000001), //i
    .io_c   (1'b0                                                                                                ), //i
    .io_s   (singleAdd_add_io_s[378:0]                                                                           ), //o
    .clk    (clk                                                                                                 ), //i
    .resetn (resetn                                                                                              )  //i
  );
  assign singleAdd_a = {_zz_singleAdd_a_20,{_zz_singleAdd_a_19,{_zz_singleAdd_a_17,{_zz_singleAdd_a_14,{_zz_singleAdd_a_10,_zz_singleAdd_a_5}}}}};
  assign io_r = _zz_io_r;
  always @(posedge clk) begin
    _zz_singleAdd_a <= io_a[63 : 0];
    _zz_singleAdd_a_1 <= _zz_singleAdd_a;
    _zz_singleAdd_a_2 <= _zz_singleAdd_a_1;
    _zz_singleAdd_a_3 <= _zz_singleAdd_a_2;
    _zz_singleAdd_a_4 <= _zz_singleAdd_a_3;
    _zz_singleAdd_a_5 <= _zz_singleAdd_a_4;
    _zz_singleAdd_a_6 <= io_a[127 : 64];
    _zz_singleAdd_a_7 <= _zz_singleAdd_a_6;
    _zz_singleAdd_a_8 <= _zz_singleAdd_a_7;
    _zz_singleAdd_a_9 <= _zz_singleAdd_a_8;
    _zz_singleAdd_a_10 <= _zz_singleAdd_a_9;
    _zz_singleAdd_a_11 <= io_a[191 : 128];
    _zz_singleAdd_a_12 <= _zz_singleAdd_a_11;
    _zz_singleAdd_a_13 <= _zz_singleAdd_a_12;
    _zz_singleAdd_a_14 <= _zz_singleAdd_a_13;
    _zz_singleAdd_a_15 <= io_a[255 : 192];
    _zz_singleAdd_a_16 <= _zz_singleAdd_a_15;
    _zz_singleAdd_a_17 <= _zz_singleAdd_a_16;
    _zz_singleAdd_a_18 <= io_a[319 : 256];
    _zz_singleAdd_a_19 <= _zz_singleAdd_a_18;
    _zz_singleAdd_a_20 <= io_a[377 : 320];
    _zz_io_r <= (singleAdd_a[377] ? _zz__zz_io_r : _zz__zz_io_r_1);
  end


endmodule

module BADD_531 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  input               io_c,
  output reg [378:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [377:0]  _zz__zz_io_s_1;
  wire       [64:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [377:0]  _zz__zz_io_s_4;
  wire       [64:0]   _zz__zz_io_s_5;
  wire       [64:0]   _zz__zz_io_s_5_1;
  wire       [0:0]    _zz__zz_io_s_5_2;
  wire       [377:0]  _zz__zz_io_s_10;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [377:0]  _zz__zz_io_s_18;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [377:0]  _zz__zz_io_s_28;
  wire       [64:0]   _zz__zz_io_s_32;
  wire       [64:0]   _zz__zz_io_s_32_1;
  wire       [0:0]    _zz__zz_io_s_32_2;
  wire       [377:0]  _zz__zz_io_s_40;
  wire       [58:0]   _zz__zz_io_s_45;
  wire       [58:0]   _zz__zz_io_s_45_1;
  wire       [0:0]    _zz__zz_io_s_45_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  wire       [64:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg        [63:0]   _zz_io_s_25;
  reg        [63:0]   _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg        [63:0]   _zz_io_s_29;
  reg        [63:0]   _zz_io_s_30;
  reg        [63:0]   _zz_io_s_31;
  wire       [64:0]   _zz_io_s_32;
  reg        [63:0]   _zz_io_s_33;
  reg                 _zz_io_s_34;
  reg        [57:0]   _zz_io_s_35;
  reg        [57:0]   _zz_io_s_36;
  reg        [57:0]   _zz_io_s_37;
  reg        [57:0]   _zz_io_s_38;
  reg        [57:0]   _zz_io_s_39;
  reg        [57:0]   _zz_io_s_40;
  reg        [57:0]   _zz_io_s_41;
  reg        [57:0]   _zz_io_s_42;
  reg        [57:0]   _zz_io_s_43;
  reg        [57:0]   _zz_io_s_44;
  wire       [58:0]   _zz_io_s_45;
  reg        [57:0]   _zz_io_s_46;
  reg                 _zz_io_s_47;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,_zz__zz_io_s_1[63 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {64'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_4 = (~ io_b);
  assign _zz__zz_io_s_5 = ({1'b0,_zz_io_s_3} + {1'b0,_zz_io_s_4});
  assign _zz__zz_io_s_5_2 = _zz_io_s_2;
  assign _zz__zz_io_s_5_1 = {64'd0, _zz__zz_io_s_5_2};
  assign _zz__zz_io_s_10 = (~ io_b);
  assign _zz__zz_io_s_12 = ({1'b0,_zz_io_s_9} + {1'b0,_zz_io_s_11});
  assign _zz__zz_io_s_12_2 = _zz_io_s_7;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_18 = (~ io_b);
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_17} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_14;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_28 = (~ io_b);
  assign _zz__zz_io_s_32 = ({1'b0,_zz_io_s_27} + {1'b0,_zz_io_s_31});
  assign _zz__zz_io_s_32_2 = _zz_io_s_23;
  assign _zz__zz_io_s_32_1 = {64'd0, _zz__zz_io_s_32_2};
  assign _zz__zz_io_s_40 = (~ io_b);
  assign _zz__zz_io_s_45 = ({1'b0,_zz_io_s_39} + {1'b0,_zz_io_s_44});
  assign _zz__zz_io_s_45_2 = _zz_io_s_34;
  assign _zz__zz_io_s_45_1 = {58'd0, _zz__zz_io_s_45_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_1;
    io_s[127 : 64] = _zz_io_s_6;
    io_s[191 : 128] = _zz_io_s_13;
    io_s[255 : 192] = _zz_io_s_22;
    io_s[319 : 256] = _zz_io_s_33;
    io_s[377 : 320] = _zz_io_s_46;
    io_s[378] = (! _zz_io_s_47);
  end

  assign _zz_io_s_5 = (_zz__zz_io_s_5 + _zz__zz_io_s_5_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_32 = (_zz__zz_io_s_32 + _zz__zz_io_s_32_1);
  assign _zz_io_s_45 = (_zz__zz_io_s_45 + _zz__zz_io_s_45_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s[64];
    _zz_io_s_3 <= io_a[127 : 64];
    _zz_io_s_4 <= _zz__zz_io_s_4[127 : 64];
    _zz_io_s_6 <= _zz_io_s_5[63:0];
    _zz_io_s_7 <= _zz_io_s_5[64];
    _zz_io_s_8 <= io_a[191 : 128];
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz__zz_io_s_10[191 : 128];
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_15 <= io_a[255 : 192];
    _zz_io_s_16 <= _zz_io_s_15;
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz__zz_io_s_18[255 : 192];
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_21[64];
    _zz_io_s_24 <= io_a[319 : 256];
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_25;
    _zz_io_s_27 <= _zz_io_s_26;
    _zz_io_s_28 <= _zz__zz_io_s_28[319 : 256];
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz_io_s_29;
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_33 <= _zz_io_s_32[63:0];
    _zz_io_s_34 <= _zz_io_s_32[64];
    _zz_io_s_35 <= io_a[377 : 320];
    _zz_io_s_36 <= _zz_io_s_35;
    _zz_io_s_37 <= _zz_io_s_36;
    _zz_io_s_38 <= _zz_io_s_37;
    _zz_io_s_39 <= _zz_io_s_38;
    _zz_io_s_40 <= _zz__zz_io_s_40[377 : 320];
    _zz_io_s_41 <= _zz_io_s_40;
    _zz_io_s_42 <= _zz_io_s_41;
    _zz_io_s_43 <= _zz_io_s_42;
    _zz_io_s_44 <= _zz_io_s_43;
    _zz_io_s_46 <= _zz_io_s_45[57:0];
    _zz_io_s_47 <= _zz_io_s_45[58];
  end


endmodule

module BADD_593 (
  input      [378:0]  io_a,
  input      [378:0]  io_b,
  input               io_c,
  output reg [379:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [378:0]  _zz__zz_io_s_1;
  wire       [64:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_8;
  wire       [378:0]  _zz__zz_io_s_8_1;
  wire       [64:0]   _zz__zz_io_s_8_2;
  wire       [0:0]    _zz__zz_io_s_8_3;
  wire       [64:0]   _zz__zz_io_s_15;
  wire       [378:0]  _zz__zz_io_s_15_1;
  wire       [64:0]   _zz__zz_io_s_15_2;
  wire       [0:0]    _zz__zz_io_s_15_3;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [378:0]  _zz__zz_io_s_21_1;
  wire       [64:0]   _zz__zz_io_s_21_2;
  wire       [0:0]    _zz__zz_io_s_21_3;
  wire       [64:0]   _zz__zz_io_s_26;
  wire       [378:0]  _zz__zz_io_s_26_1;
  wire       [64:0]   _zz__zz_io_s_26_2;
  wire       [0:0]    _zz__zz_io_s_26_3;
  wire       [59:0]   _zz__zz_io_s_30;
  wire       [378:0]  _zz__zz_io_s_30_1;
  wire       [59:0]   _zz__zz_io_s_30_2;
  wire       [0:0]    _zz__zz_io_s_30_3;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  wire       [64:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [64:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg                 _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg        [63:0]   _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg                 _zz_io_s_25;
  wire       [64:0]   _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg                 _zz_io_s_29;
  wire       [59:0]   _zz_io_s_30;
  reg        [58:0]   _zz_io_s_31;
  reg                 _zz_io_s_32;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,_zz__zz_io_s_1[63 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {64'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_8 = ({1'b0,io_a[127 : 64]} + {1'b0,_zz__zz_io_s_8_1[127 : 64]});
  assign _zz__zz_io_s_8_1 = (~ io_b);
  assign _zz__zz_io_s_8_3 = _zz_io_s_7;
  assign _zz__zz_io_s_8_2 = {64'd0, _zz__zz_io_s_8_3};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[191 : 128]} + {1'b0,_zz__zz_io_s_15_1[191 : 128]});
  assign _zz__zz_io_s_15_1 = (~ io_b);
  assign _zz__zz_io_s_15_3 = _zz_io_s_14;
  assign _zz__zz_io_s_15_2 = {64'd0, _zz__zz_io_s_15_3};
  assign _zz__zz_io_s_21 = ({1'b0,io_a[255 : 192]} + {1'b0,_zz__zz_io_s_21_1[255 : 192]});
  assign _zz__zz_io_s_21_1 = (~ io_b);
  assign _zz__zz_io_s_21_3 = _zz_io_s_20;
  assign _zz__zz_io_s_21_2 = {64'd0, _zz__zz_io_s_21_3};
  assign _zz__zz_io_s_26 = ({1'b0,io_a[319 : 256]} + {1'b0,_zz__zz_io_s_26_1[319 : 256]});
  assign _zz__zz_io_s_26_1 = (~ io_b);
  assign _zz__zz_io_s_26_3 = _zz_io_s_25;
  assign _zz__zz_io_s_26_2 = {64'd0, _zz__zz_io_s_26_3};
  assign _zz__zz_io_s_30 = ({1'b0,io_a[378 : 320]} + {1'b0,_zz__zz_io_s_30_1[378 : 320]});
  assign _zz__zz_io_s_30_1 = (~ io_b);
  assign _zz__zz_io_s_30_3 = _zz_io_s_29;
  assign _zz__zz_io_s_30_2 = {59'd0, _zz__zz_io_s_30_3};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_6;
    io_s[127 : 64] = _zz_io_s_13;
    io_s[191 : 128] = _zz_io_s_19;
    io_s[255 : 192] = _zz_io_s_24;
    io_s[319 : 256] = _zz_io_s_28;
    io_s[378 : 320] = _zz_io_s_31;
    io_s[379] = (! _zz_io_s_32);
  end

  assign _zz_io_s_8 = (_zz__zz_io_s_8 + _zz__zz_io_s_8_2);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_2);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_2);
  assign _zz_io_s_26 = (_zz__zz_io_s_26 + _zz__zz_io_s_26_2);
  assign _zz_io_s_30 = (_zz__zz_io_s_30 + _zz__zz_io_s_30_2);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= _zz_io_s[64];
    _zz_io_s_9 <= _zz_io_s_8[63:0];
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= _zz_io_s_11;
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_8[64];
    _zz_io_s_16 <= _zz_io_s_15[63:0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_15[64];
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_22;
    _zz_io_s_24 <= _zz_io_s_23;
    _zz_io_s_25 <= _zz_io_s_21[64];
    _zz_io_s_27 <= _zz_io_s_26[63:0];
    _zz_io_s_28 <= _zz_io_s_27;
    _zz_io_s_29 <= _zz_io_s_26[64];
    _zz_io_s_31 <= _zz_io_s_30[58:0];
    _zz_io_s_32 <= _zz_io_s_30[59];
  end


endmodule

module BADD_592 (
  input      [120:0]  io_a,
  input      [120:0]  io_b,
  input               io_c,
  output reg [121:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [62:0]   _zz__zz_io_s;
  wire       [62:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [62:0]   _zz_io_s;
  reg        [61:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[61 : 0]} + {1'b0,io_b[61 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {62'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[120 : 62]} + {1'b0,io_b[120 : 62]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[61 : 0] = _zz_io_s_1;
    io_s[120 : 62] = _zz_io_s_4;
    io_s[121] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[61:0];
    _zz_io_s_2 <= _zz_io_s[62];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_591 (
  input      [36:0]   io_a,
  input      [36:0]   io_b,
  input               io_c,
  output reg [37:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [37:0]   _zz__zz_io_s;
  wire       [37:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [37:0]   _zz_io_s;
  reg        [36:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[36 : 0]} + {1'b0,io_b[36 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {37'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[36 : 0] = _zz_io_s_1;
    io_s[37] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[36:0];
    _zz_io_s_2 <= _zz_io_s[37];
  end


endmodule

module BADD_590 (
  input      [9:0]    io_a,
  input      [9:0]    io_b,
  input               io_c,
  output reg [10:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [10:0]   _zz__zz_io_s;
  wire       [10:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [10:0]   _zz_io_s;
  reg        [9:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[9 : 0]} + {1'b0,io_b[9 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {10'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[9 : 0] = _zz_io_s_1;
    io_s[10] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[9:0];
    _zz_io_s_2 <= _zz_io_s[10];
  end


endmodule

module BADD_589 (
  input      [68:0]   io_a,
  input      [68:0]   io_b,
  input               io_c,
  output reg [69:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [10:0]   _zz__zz_io_s;
  wire       [10:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [10:0]   _zz_io_s;
  reg        [9:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[9 : 0]} + {1'b0,io_b[9 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {10'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[68 : 10]} + {1'b0,io_b[68 : 10]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[9 : 0] = _zz_io_s_1;
    io_s[68 : 10] = _zz_io_s_4;
    io_s[69] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[9:0];
    _zz_io_s_2 <= _zz_io_s[10];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_588 (
  input      [58:0]   io_a,
  input      [58:0]   io_b,
  input               io_c,
  output reg [59:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [59:0]   _zz__zz_io_s;
  wire       [59:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz_io_s;
  reg        [58:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[58 : 0]} + {1'b0,io_b[58 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {59'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[58 : 0] = _zz_io_s_1;
    io_s[59] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[58:0];
    _zz_io_s_2 <= _zz_io_s[59];
  end


endmodule

module BADD_587 (
  input      [54:0]   io_a,
  input      [54:0]   io_b,
  input               io_c,
  output reg [55:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [55:0]   _zz__zz_io_s;
  wire       [55:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [55:0]   _zz_io_s;
  reg        [54:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[54 : 0]} + {1'b0,io_b[54 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {55'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[54 : 0] = _zz_io_s_1;
    io_s[55] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[54:0];
    _zz_io_s_2 <= _zz_io_s[55];
  end


endmodule

module BADD_586 (
  input      [63:0]   io_a,
  input      [63:0]   io_b,
  input               io_c,
  output reg [64:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [5:0]    _zz__zz_io_s;
  wire       [5:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [5:0]    _zz_io_s;
  reg        [4:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[4 : 0]} + {1'b0,io_b[4 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {5'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[63 : 5]} + {1'b0,io_b[63 : 5]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[4 : 0] = _zz_io_s_1;
    io_s[63 : 5] = _zz_io_s_4;
    io_s[64] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[4:0];
    _zz_io_s_2 <= _zz_io_s[5];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_585 (
  input      [84:0]   io_a,
  input      [84:0]   io_b,
  input               io_c,
  output reg [85:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [26:0]   _zz__zz_io_s;
  wire       [26:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [26:0]   _zz_io_s;
  reg        [25:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[25 : 0]} + {1'b0,io_b[25 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {26'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[84 : 26]} + {1'b0,io_b[84 : 26]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[25 : 0] = _zz_io_s_1;
    io_s[84 : 26] = _zz_io_s_4;
    io_s[85] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[25:0];
    _zz_io_s_2 <= _zz_io_s[26];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_584 (
  input      [74:0]   io_a,
  input      [74:0]   io_b,
  input               io_c,
  output reg [75:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [16:0]   _zz__zz_io_s;
  wire       [16:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [16:0]   _zz_io_s;
  reg        [15:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[15 : 0]} + {1'b0,io_b[15 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {16'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[74 : 16]} + {1'b0,io_b[74 : 16]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[15 : 0] = _zz_io_s_1;
    io_s[74 : 16] = _zz_io_s_4;
    io_s[75] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[15:0];
    _zz_io_s_2 <= _zz_io_s[16];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_583 (
  input      [96:0]   io_a,
  input      [96:0]   io_b,
  input               io_c,
  output reg [97:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [38:0]   _zz__zz_io_s;
  wire       [38:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [38:0]   _zz_io_s;
  reg        [37:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[37 : 0]} + {1'b0,io_b[37 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {38'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[96 : 38]} + {1'b0,io_b[96 : 38]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[37 : 0] = _zz_io_s_1;
    io_s[96 : 38] = _zz_io_s_4;
    io_s[97] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[37:0];
    _zz_io_s_2 <= _zz_io_s[38];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_582 (
  input      [189:0]  io_a,
  input      [189:0]  io_b,
  input               io_c,
  output reg [190:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [3:0]    _zz__zz_io_s;
  wire       [3:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [3:0]    _zz_io_s;
  reg        [2:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[2 : 0]} + {1'b0,io_b[2 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {3'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[66 : 3]} + {1'b0,io_b[66 : 3]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[130 : 67]} + {1'b0,io_b[130 : 67]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[189 : 131]} + {1'b0,io_b[189 : 131]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[2 : 0] = _zz_io_s_1;
    io_s[66 : 3] = _zz_io_s_4;
    io_s[130 : 67] = _zz_io_s_7;
    io_s[189 : 131] = _zz_io_s_10;
    io_s[190] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[2:0];
    _zz_io_s_2 <= _zz_io_s[3];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_581 (
  input      [145:0]  io_a,
  input      [145:0]  io_b,
  input               io_c,
  output reg [146:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [23:0]   _zz__zz_io_s;
  wire       [23:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [23:0]   _zz_io_s;
  reg        [22:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[22 : 0]} + {1'b0,io_b[22 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {23'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[86 : 23]} + {1'b0,io_b[86 : 23]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[145 : 87]} + {1'b0,io_b[145 : 87]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[22 : 0] = _zz_io_s_1;
    io_s[86 : 23] = _zz_io_s_4;
    io_s[145 : 87] = _zz_io_s_7;
    io_s[146] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[22:0];
    _zz_io_s_2 <= _zz_io_s[23];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_580 (
  input      [129:0]  io_a,
  input      [129:0]  io_b,
  input               io_c,
  output reg [130:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [7:0]    _zz__zz_io_s;
  wire       [7:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [7:0]    _zz_io_s;
  reg        [6:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[6 : 0]} + {1'b0,io_b[6 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {7'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[70 : 7]} + {1'b0,io_b[70 : 7]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[129 : 71]} + {1'b0,io_b[129 : 71]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[6 : 0] = _zz_io_s_1;
    io_s[70 : 7] = _zz_io_s_4;
    io_s[129 : 71] = _zz_io_s_7;
    io_s[130] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[6:0];
    _zz_io_s_2 <= _zz_io_s[7];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_579 (
  input      [125:0]  io_a,
  input      [125:0]  io_b,
  input               io_c,
  output reg [126:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [3:0]    _zz__zz_io_s;
  wire       [3:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [3:0]    _zz_io_s;
  reg        [2:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[2 : 0]} + {1'b0,io_b[2 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {3'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[66 : 3]} + {1'b0,io_b[66 : 3]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[125 : 67]} + {1'b0,io_b[125 : 67]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[2 : 0] = _zz_io_s_1;
    io_s[66 : 3] = _zz_io_s_4;
    io_s[125 : 67] = _zz_io_s_7;
    io_s[126] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[2:0];
    _zz_io_s_2 <= _zz_io_s[3];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_578 (
  input      [141:0]  io_a,
  input      [141:0]  io_b,
  input               io_c,
  output reg [142:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [19:0]   _zz__zz_io_s;
  wire       [19:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [19:0]   _zz_io_s;
  reg        [18:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[18 : 0]} + {1'b0,io_b[18 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {19'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[82 : 19]} + {1'b0,io_b[82 : 19]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[141 : 83]} + {1'b0,io_b[141 : 83]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[18 : 0] = _zz_io_s_1;
    io_s[82 : 19] = _zz_io_s_4;
    io_s[141 : 83] = _zz_io_s_7;
    io_s[142] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[18:0];
    _zz_io_s_2 <= _zz_io_s[19];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_577 (
  input      [166:0]  io_a,
  input      [166:0]  io_b,
  input               io_c,
  output reg [167:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [44:0]   _zz__zz_io_s;
  wire       [44:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [44:0]   _zz_io_s;
  reg        [43:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[43 : 0]} + {1'b0,io_b[43 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {44'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[107 : 44]} + {1'b0,io_b[107 : 44]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[166 : 108]} + {1'b0,io_b[166 : 108]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[43 : 0] = _zz_io_s_1;
    io_s[107 : 44] = _zz_io_s_4;
    io_s[166 : 108] = _zz_io_s_7;
    io_s[167] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[43:0];
    _zz_io_s_2 <= _zz_io_s[44];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_576 (
  input      [150:0]  io_a,
  input      [150:0]  io_b,
  input               io_c,
  output reg [151:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [28:0]   _zz__zz_io_s;
  wire       [28:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [28:0]   _zz_io_s;
  reg        [27:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[27 : 0]} + {1'b0,io_b[27 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {28'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[91 : 28]} + {1'b0,io_b[91 : 28]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[150 : 92]} + {1'b0,io_b[150 : 92]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[27 : 0] = _zz_io_s_1;
    io_s[91 : 28] = _zz_io_s_4;
    io_s[150 : 92] = _zz_io_s_7;
    io_s[151] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[27:0];
    _zz_io_s_2 <= _zz_io_s[28];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_575 (
  input      [182:0]  io_a,
  input      [182:0]  io_b,
  input               io_c,
  output reg [183:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [60:0]   _zz__zz_io_s;
  wire       [60:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [60:0]   _zz_io_s;
  reg        [59:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[59 : 0]} + {1'b0,io_b[59 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {60'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[123 : 60]} + {1'b0,io_b[123 : 60]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[182 : 124]} + {1'b0,io_b[182 : 124]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[59 : 0] = _zz_io_s_1;
    io_s[123 : 60] = _zz_io_s_4;
    io_s[182 : 124] = _zz_io_s_7;
    io_s[183] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[59:0];
    _zz_io_s_2 <= _zz_io_s[60];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_574 (
  input      [220:0]  io_a,
  input      [220:0]  io_b,
  input               io_c,
  output reg [221:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [34:0]   _zz__zz_io_s;
  wire       [34:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [34:0]   _zz_io_s;
  reg        [33:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[33 : 0]} + {1'b0,io_b[33 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {34'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[97 : 34]} + {1'b0,io_b[97 : 34]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[161 : 98]} + {1'b0,io_b[161 : 98]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[220 : 162]} + {1'b0,io_b[220 : 162]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[33 : 0] = _zz_io_s_1;
    io_s[97 : 34] = _zz_io_s_4;
    io_s[161 : 98] = _zz_io_s_7;
    io_s[220 : 162] = _zz_io_s_10;
    io_s[221] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[33:0];
    _zz_io_s_2 <= _zz_io_s[34];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_573 (
  input      [200:0]  io_a,
  input      [200:0]  io_b,
  input               io_c,
  output reg [201:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [14:0]   _zz__zz_io_s;
  wire       [14:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [14:0]   _zz_io_s;
  reg        [13:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[13 : 0]} + {1'b0,io_b[13 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {14'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[77 : 14]} + {1'b0,io_b[77 : 14]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[141 : 78]} + {1'b0,io_b[141 : 78]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[200 : 142]} + {1'b0,io_b[200 : 142]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[13 : 0] = _zz_io_s_1;
    io_s[77 : 14] = _zz_io_s_4;
    io_s[141 : 78] = _zz_io_s_7;
    io_s[200 : 142] = _zz_io_s_10;
    io_s[201] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[13:0];
    _zz_io_s_2 <= _zz_io_s[14];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_572 (
  input      [194:0]  io_a,
  input      [194:0]  io_b,
  input               io_c,
  output reg [195:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [8:0]    _zz__zz_io_s;
  wire       [8:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [8:0]    _zz_io_s;
  reg        [7:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[7 : 0]} + {1'b0,io_b[7 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {8'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[71 : 8]} + {1'b0,io_b[71 : 8]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[135 : 72]} + {1'b0,io_b[135 : 72]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[194 : 136]} + {1'b0,io_b[194 : 136]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[7 : 0] = _zz_io_s_1;
    io_s[71 : 8] = _zz_io_s_4;
    io_s[135 : 72] = _zz_io_s_7;
    io_s[194 : 136] = _zz_io_s_10;
    io_s[195] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[7:0];
    _zz_io_s_2 <= _zz_io_s[8];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_571 (
  input      [205:0]  io_a,
  input      [205:0]  io_b,
  input               io_c,
  output reg [206:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [19:0]   _zz__zz_io_s;
  wire       [19:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [19:0]   _zz_io_s;
  reg        [18:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[18 : 0]} + {1'b0,io_b[18 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {19'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[82 : 19]} + {1'b0,io_b[82 : 19]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[146 : 83]} + {1'b0,io_b[146 : 83]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[205 : 147]} + {1'b0,io_b[205 : 147]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[18 : 0] = _zz_io_s_1;
    io_s[82 : 19] = _zz_io_s_4;
    io_s[146 : 83] = _zz_io_s_7;
    io_s[205 : 147] = _zz_io_s_10;
    io_s[206] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[18:0];
    _zz_io_s_2 <= _zz_io_s[19];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_570 (
  input      [258:0]  io_a,
  input      [258:0]  io_b,
  input               io_c,
  output reg [259:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [8:0]    _zz__zz_io_s;
  wire       [8:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [59:0]   _zz__zz_io_s_12;
  wire       [59:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [8:0]    _zz_io_s;
  reg        [7:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [59:0]   _zz_io_s_12;
  reg        [58:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[7 : 0]} + {1'b0,io_b[7 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {8'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[71 : 8]} + {1'b0,io_b[71 : 8]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[135 : 72]} + {1'b0,io_b[135 : 72]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[199 : 136]} + {1'b0,io_b[199 : 136]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[258 : 200]} + {1'b0,io_b[258 : 200]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {59'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[7 : 0] = _zz_io_s_1;
    io_s[71 : 8] = _zz_io_s_4;
    io_s[135 : 72] = _zz_io_s_7;
    io_s[199 : 136] = _zz_io_s_10;
    io_s[258 : 200] = _zz_io_s_13;
    io_s[259] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[7:0];
    _zz_io_s_2 <= _zz_io_s[8];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[58:0];
    _zz_io_s_14 <= _zz_io_s_12[59];
  end


endmodule

module BADD_569 (
  input      [225:0]  io_a,
  input      [225:0]  io_b,
  input               io_c,
  output reg [226:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [39:0]   _zz__zz_io_s;
  wire       [39:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [39:0]   _zz_io_s;
  reg        [38:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[38 : 0]} + {1'b0,io_b[38 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {39'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[102 : 39]} + {1'b0,io_b[102 : 39]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[166 : 103]} + {1'b0,io_b[166 : 103]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[225 : 167]} + {1'b0,io_b[225 : 167]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[38 : 0] = _zz_io_s_1;
    io_s[102 : 39] = _zz_io_s_4;
    io_s[166 : 103] = _zz_io_s_7;
    io_s[225 : 167] = _zz_io_s_10;
    io_s[226] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[38:0];
    _zz_io_s_2 <= _zz_io_s[39];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_568 (
  input      [267:0]  io_a,
  input      [267:0]  io_b,
  input               io_c,
  output reg [268:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [17:0]   _zz__zz_io_s;
  wire       [17:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [59:0]   _zz__zz_io_s_12;
  wire       [59:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [17:0]   _zz_io_s;
  reg        [16:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [59:0]   _zz_io_s_12;
  reg        [58:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[16 : 0]} + {1'b0,io_b[16 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {17'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[80 : 17]} + {1'b0,io_b[80 : 17]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[144 : 81]} + {1'b0,io_b[144 : 81]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[208 : 145]} + {1'b0,io_b[208 : 145]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[267 : 209]} + {1'b0,io_b[267 : 209]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {59'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[16 : 0] = _zz_io_s_1;
    io_s[80 : 17] = _zz_io_s_4;
    io_s[144 : 81] = _zz_io_s_7;
    io_s[208 : 145] = _zz_io_s_10;
    io_s[267 : 209] = _zz_io_s_13;
    io_s[268] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[16:0];
    _zz_io_s_2 <= _zz_io_s[17];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[58:0];
    _zz_io_s_14 <= _zz_io_s_12[59];
  end


endmodule

module BADD_567 (
  input      [4:0]    io_a,
  input      [4:0]    io_b,
  input               io_c,
  output reg [5:0]    io_s,
  input               clk,
  input               resetn
);

  wire       [5:0]    _zz__zz_io_s;
  wire       [5:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [5:0]    _zz_io_s;
  reg        [4:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[4 : 0]} + {1'b0,io_b[4 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {5'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[4 : 0] = _zz_io_s_1;
    io_s[5] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[4:0];
    _zz_io_s_2 <= _zz_io_s[5];
  end


endmodule

module BADD_566 (
  input      [162:0]  io_a,
  input      [162:0]  io_b,
  input               io_c,
  output reg [163:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [40:0]   _zz__zz_io_s;
  wire       [40:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [40:0]   _zz_io_s;
  reg        [39:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[39 : 0]} + {1'b0,io_b[39 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {40'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[103 : 40]} + {1'b0,io_b[103 : 40]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[162 : 104]} + {1'b0,io_b[162 : 104]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[39 : 0] = _zz_io_s_1;
    io_s[103 : 40] = _zz_io_s_4;
    io_s[162 : 104] = _zz_io_s_7;
    io_s[163] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[39:0];
    _zz_io_s_2 <= _zz_io_s[40];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_565 (
  input      [79:0]   io_a,
  input      [79:0]   io_b,
  input               io_c,
  output reg [80:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [21:0]   _zz__zz_io_s;
  wire       [21:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [21:0]   _zz_io_s;
  reg        [20:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[20 : 0]} + {1'b0,io_b[20 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {21'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[79 : 21]} + {1'b0,io_b[79 : 21]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[20 : 0] = _zz_io_s_1;
    io_s[79 : 21] = _zz_io_s_4;
    io_s[80] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[20:0];
    _zz_io_s_2 <= _zz_io_s[21];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_564 (
  input      [31:0]   io_a,
  input      [31:0]   io_b,
  input               io_c,
  output reg [32:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [32:0]   _zz__zz_io_s;
  wire       [32:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [32:0]   _zz_io_s;
  reg        [31:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[31 : 0]} + {1'b0,io_b[31 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {32'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[31 : 0] = _zz_io_s_1;
    io_s[32] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[31:0];
    _zz_io_s_2 <= _zz_io_s[32];
  end


endmodule

module BADD_563 (
  input      [20:0]   io_a,
  input      [20:0]   io_b,
  input               io_c,
  output reg [21:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [21:0]   _zz__zz_io_s;
  wire       [21:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [21:0]   _zz_io_s;
  reg        [20:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[20 : 0]} + {1'b0,io_b[20 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {21'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[20 : 0] = _zz_io_s_1;
    io_s[21] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[20:0];
    _zz_io_s_2 <= _zz_io_s[21];
  end


endmodule

module BADD_562 (
  input      [15:0]   io_a,
  input      [15:0]   io_b,
  input               io_c,
  output reg [16:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [16:0]   _zz__zz_io_s;
  wire       [16:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [16:0]   _zz_io_s;
  reg        [15:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[15 : 0]} + {1'b0,io_b[15 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {16'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[15 : 0] = _zz_io_s_1;
    io_s[16] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[15:0];
    _zz_io_s_2 <= _zz_io_s[16];
  end


endmodule

module BADD_561 (
  input      [25:0]   io_a,
  input      [25:0]   io_b,
  input               io_c,
  output reg [26:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [26:0]   _zz__zz_io_s;
  wire       [26:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [26:0]   _zz_io_s;
  reg        [25:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[25 : 0]} + {1'b0,io_b[25 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {26'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[25 : 0] = _zz_io_s_1;
    io_s[26] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[25:0];
    _zz_io_s_2 <= _zz_io_s[26];
  end


endmodule

module BADD_560 (
  input      [46:0]   io_a,
  input      [46:0]   io_b,
  input               io_c,
  output reg [47:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [47:0]   _zz__zz_io_s;
  wire       [47:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [47:0]   _zz_io_s;
  reg        [46:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[46 : 0]} + {1'b0,io_b[46 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {47'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[46 : 0] = _zz_io_s_1;
    io_s[47] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[46:0];
    _zz_io_s_2 <= _zz_io_s[47];
  end


endmodule

module BADD_559 (
  input      [42:0]   io_a,
  input      [42:0]   io_b,
  input               io_c,
  output reg [43:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [43:0]   _zz__zz_io_s;
  wire       [43:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [43:0]   _zz_io_s;
  reg        [42:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[42 : 0]} + {1'b0,io_b[42 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {43'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[42 : 0] = _zz_io_s_1;
    io_s[43] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[42:0];
    _zz_io_s_2 <= _zz_io_s[43];
  end


endmodule

module BADD_558 (
  input      [50:0]   io_a,
  input      [50:0]   io_b,
  input               io_c,
  output reg [51:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [51:0]   _zz__zz_io_s;
  wire       [51:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [51:0]   _zz_io_s;
  reg        [50:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;

  assign _zz__zz_io_s = ({1'b0,io_a[50 : 0]} + {1'b0,io_b[50 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {51'd0, _zz__zz_io_s_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[50 : 0] = _zz_io_s_1;
    io_s[51] = _zz_io_s_2;
  end

  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[50:0];
    _zz_io_s_2 <= _zz_io_s[51];
  end


endmodule

module BADD_557 (
  input      [111:0]  io_a,
  input      [111:0]  io_b,
  input               io_c,
  output reg [112:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [53:0]   _zz__zz_io_s;
  wire       [53:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [53:0]   _zz_io_s;
  reg        [52:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[52 : 0]} + {1'b0,io_b[52 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {53'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[111 : 53]} + {1'b0,io_b[111 : 53]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[52 : 0] = _zz_io_s_1;
    io_s[111 : 53] = _zz_io_s_4;
    io_s[112] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[52:0];
    _zz_io_s_2 <= _zz_io_s[53];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_556 (
  input      [101:0]  io_a,
  input      [101:0]  io_b,
  input               io_c,
  output reg [102:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [43:0]   _zz__zz_io_s;
  wire       [43:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [43:0]   _zz_io_s;
  reg        [42:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[42 : 0]} + {1'b0,io_b[42 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {43'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[101 : 43]} + {1'b0,io_b[101 : 43]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[42 : 0] = _zz_io_s_1;
    io_s[101 : 43] = _zz_io_s_4;
    io_s[102] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[42:0];
    _zz_io_s_2 <= _zz_io_s[43];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_555 (
  input      [91:0]   io_a,
  input      [91:0]   io_b,
  input               io_c,
  output reg [92:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [33:0]   _zz__zz_io_s;
  wire       [33:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [33:0]   _zz_io_s;
  reg        [32:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[32 : 0]} + {1'b0,io_b[32 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {33'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[91 : 33]} + {1'b0,io_b[91 : 33]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[32 : 0] = _zz_io_s_1;
    io_s[91 : 33] = _zz_io_s_4;
    io_s[92] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[32:0];
    _zz_io_s_2 <= _zz_io_s[33];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_554 (
  input      [106:0]  io_a,
  input      [106:0]  io_b,
  input               io_c,
  output reg [107:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[106 : 48]} + {1'b0,io_b[106 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[106 : 48] = _zz_io_s_4;
    io_s[107] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_553 (
  input      [136:0]  io_a,
  input      [136:0]  io_b,
  input               io_c,
  output reg [137:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [14:0]   _zz__zz_io_s;
  wire       [14:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [14:0]   _zz_io_s;
  reg        [13:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[13 : 0]} + {1'b0,io_b[13 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {14'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[77 : 14]} + {1'b0,io_b[77 : 14]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[136 : 78]} + {1'b0,io_b[136 : 78]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[13 : 0] = _zz_io_s_1;
    io_s[77 : 14] = _zz_io_s_4;
    io_s[136 : 78] = _zz_io_s_7;
    io_s[137] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[13:0];
    _zz_io_s_2 <= _zz_io_s[14];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_552 (
  input      [116:0]  io_a,
  input      [116:0]  io_b,
  input               io_c,
  output reg [117:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [58:0]   _zz__zz_io_s;
  wire       [58:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [59:0]   _zz__zz_io_s_3;
  wire       [59:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [58:0]   _zz_io_s;
  reg        [57:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [59:0]   _zz_io_s_3;
  reg        [58:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;

  assign _zz__zz_io_s = ({1'b0,io_a[57 : 0]} + {1'b0,io_b[57 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {58'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[116 : 58]} + {1'b0,io_b[116 : 58]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {59'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[57 : 0] = _zz_io_s_1;
    io_s[116 : 58] = _zz_io_s_4;
    io_s[117] = _zz_io_s_5;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[57:0];
    _zz_io_s_2 <= _zz_io_s[58];
    _zz_io_s_4 <= _zz_io_s_3[58:0];
    _zz_io_s_5 <= _zz_io_s_3[59];
  end


endmodule

module BADD_551 (
  input      [154:0]  io_a,
  input      [154:0]  io_b,
  input               io_c,
  output reg [155:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [32:0]   _zz__zz_io_s;
  wire       [32:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [32:0]   _zz_io_s;
  reg        [31:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[31 : 0]} + {1'b0,io_b[31 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {32'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 32]} + {1'b0,io_b[95 : 32]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[154 : 96]} + {1'b0,io_b[154 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[31 : 0] = _zz_io_s_1;
    io_s[95 : 32] = _zz_io_s_4;
    io_s[154 : 96] = _zz_io_s_7;
    io_s[155] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[31:0];
    _zz_io_s_2 <= _zz_io_s[32];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_550 (
  input      [262:0]  io_a,
  input      [262:0]  io_b,
  input               io_c,
  output reg [263:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [12:0]   _zz__zz_io_s;
  wire       [12:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [59:0]   _zz__zz_io_s_12;
  wire       [59:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [12:0]   _zz_io_s;
  reg        [11:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [59:0]   _zz_io_s_12;
  reg        [58:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[11 : 0]} + {1'b0,io_b[11 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {12'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[75 : 12]} + {1'b0,io_b[75 : 12]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[139 : 76]} + {1'b0,io_b[139 : 76]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[203 : 140]} + {1'b0,io_b[203 : 140]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[262 : 204]} + {1'b0,io_b[262 : 204]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {59'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[11 : 0] = _zz_io_s_1;
    io_s[75 : 12] = _zz_io_s_4;
    io_s[139 : 76] = _zz_io_s_7;
    io_s[203 : 140] = _zz_io_s_10;
    io_s[262 : 204] = _zz_io_s_13;
    io_s[263] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[11:0];
    _zz_io_s_2 <= _zz_io_s[12];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[58:0];
    _zz_io_s_14 <= _zz_io_s_12[59];
  end


endmodule

module BADD_549 (
  input      [214:0]  io_a,
  input      [214:0]  io_b,
  input               io_c,
  output reg [215:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [28:0]   _zz__zz_io_s;
  wire       [28:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [28:0]   _zz_io_s;
  reg        [27:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[27 : 0]} + {1'b0,io_b[27 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {28'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[91 : 28]} + {1'b0,io_b[91 : 28]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[155 : 92]} + {1'b0,io_b[155 : 92]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[214 : 156]} + {1'b0,io_b[214 : 156]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[27 : 0] = _zz_io_s_1;
    io_s[91 : 28] = _zz_io_s_4;
    io_s[155 : 92] = _zz_io_s_7;
    io_s[214 : 156] = _zz_io_s_10;
    io_s[215] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[27:0];
    _zz_io_s_2 <= _zz_io_s[28];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_548 (
  input      [176:0]  io_a,
  input      [176:0]  io_b,
  input               io_c,
  output reg [177:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [54:0]   _zz__zz_io_s;
  wire       [54:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [54:0]   _zz_io_s;
  reg        [53:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[53 : 0]} + {1'b0,io_b[53 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {54'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[117 : 54]} + {1'b0,io_b[117 : 54]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[176 : 118]} + {1'b0,io_b[176 : 118]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[53 : 0] = _zz_io_s_1;
    io_s[117 : 54] = _zz_io_s_4;
    io_s[176 : 118] = _zz_io_s_7;
    io_s[177] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[53:0];
    _zz_io_s_2 <= _zz_io_s[54];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_547 (
  input      [170:0]  io_a,
  input      [170:0]  io_b,
  input               io_c,
  output reg [171:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [59:0]   _zz__zz_io_s_6;
  wire       [59:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [59:0]   _zz_io_s_6;
  reg        [58:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[111 : 48]} + {1'b0,io_b[111 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[170 : 112]} + {1'b0,io_b[170 : 112]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {59'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[111 : 48] = _zz_io_s_4;
    io_s[170 : 112] = _zz_io_s_7;
    io_s[171] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[58:0];
    _zz_io_s_8 <= _zz_io_s_6[59];
  end


endmodule

module BADD_546 (
  input      [209:0]  io_a,
  input      [209:0]  io_b,
  input               io_c,
  output reg [210:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [23:0]   _zz__zz_io_s;
  wire       [23:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [23:0]   _zz_io_s;
  reg        [22:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[22 : 0]} + {1'b0,io_b[22 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {23'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[86 : 23]} + {1'b0,io_b[86 : 23]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[150 : 87]} + {1'b0,io_b[150 : 87]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[209 : 151]} + {1'b0,io_b[209 : 151]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[22 : 0] = _zz_io_s_1;
    io_s[86 : 23] = _zz_io_s_4;
    io_s[150 : 87] = _zz_io_s_7;
    io_s[209 : 151] = _zz_io_s_10;
    io_s[210] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[22:0];
    _zz_io_s_2 <= _zz_io_s[23];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_545 (
  input      [239:0]  io_a,
  input      [239:0]  io_b,
  input               io_c,
  output reg [240:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [53:0]   _zz__zz_io_s;
  wire       [53:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [53:0]   _zz_io_s;
  reg        [52:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[52 : 0]} + {1'b0,io_b[52 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {53'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[116 : 53]} + {1'b0,io_b[116 : 53]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[180 : 117]} + {1'b0,io_b[180 : 117]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[239 : 181]} + {1'b0,io_b[239 : 181]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[52 : 0] = _zz_io_s_1;
    io_s[116 : 53] = _zz_io_s_4;
    io_s[180 : 117] = _zz_io_s_7;
    io_s[239 : 181] = _zz_io_s_10;
    io_s[240] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[52:0];
    _zz_io_s_2 <= _zz_io_s[53];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_544 (
  input      [234:0]  io_a,
  input      [234:0]  io_b,
  input               io_c,
  output reg [235:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [59:0]   _zz__zz_io_s_9;
  wire       [59:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [59:0]   _zz_io_s_9;
  reg        [58:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[111 : 48]} + {1'b0,io_b[111 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[175 : 112]} + {1'b0,io_b[175 : 112]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[234 : 176]} + {1'b0,io_b[234 : 176]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {59'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[111 : 48] = _zz_io_s_4;
    io_s[175 : 112] = _zz_io_s_7;
    io_s[234 : 176] = _zz_io_s_10;
    io_s[235] = _zz_io_s_11;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[58:0];
    _zz_io_s_11 <= _zz_io_s_9[59];
  end


endmodule

module BADD_543 (
  input      [253:0]  io_a,
  input      [253:0]  io_b,
  input               io_c,
  output reg [254:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [3:0]    _zz__zz_io_s;
  wire       [3:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [59:0]   _zz__zz_io_s_12;
  wire       [59:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [3:0]    _zz_io_s;
  reg        [2:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [59:0]   _zz_io_s_12;
  reg        [58:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[2 : 0]} + {1'b0,io_b[2 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {3'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[66 : 3]} + {1'b0,io_b[66 : 3]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[130 : 67]} + {1'b0,io_b[130 : 67]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[194 : 131]} + {1'b0,io_b[194 : 131]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[253 : 195]} + {1'b0,io_b[253 : 195]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {59'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[2 : 0] = _zz_io_s_1;
    io_s[66 : 3] = _zz_io_s_4;
    io_s[130 : 67] = _zz_io_s_7;
    io_s[194 : 131] = _zz_io_s_10;
    io_s[253 : 195] = _zz_io_s_13;
    io_s[254] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[2:0];
    _zz_io_s_2 <= _zz_io_s[3];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[58:0];
    _zz_io_s_14 <= _zz_io_s_12[59];
  end


endmodule

module BADD_542 (
  input      [315:0]  io_a,
  input      [315:0]  io_b,
  input               io_c,
  output reg [316:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [1:0]    _zz__zz_io_s;
  wire       [1:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [59:0]   _zz__zz_io_s_15;
  wire       [59:0]   _zz__zz_io_s_15_1;
  wire       [0:0]    _zz__zz_io_s_15_2;
  wire       [1:0]    _zz_io_s;
  reg        [0:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [59:0]   _zz_io_s_15;
  reg        [58:0]   _zz_io_s_16;
  reg                 _zz_io_s_17;

  assign _zz__zz_io_s = ({1'b0,io_a[0 : 0]} + {1'b0,io_b[0 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {1'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[64 : 1]} + {1'b0,io_b[64 : 1]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[128 : 65]} + {1'b0,io_b[128 : 65]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[192 : 129]} + {1'b0,io_b[192 : 129]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[256 : 193]} + {1'b0,io_b[256 : 193]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[315 : 257]} + {1'b0,io_b[315 : 257]});
  assign _zz__zz_io_s_15_2 = _zz_io_s_14;
  assign _zz__zz_io_s_15_1 = {59'd0, _zz__zz_io_s_15_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[0 : 0] = _zz_io_s_1;
    io_s[64 : 1] = _zz_io_s_4;
    io_s[128 : 65] = _zz_io_s_7;
    io_s[192 : 129] = _zz_io_s_10;
    io_s[256 : 193] = _zz_io_s_13;
    io_s[315 : 257] = _zz_io_s_16;
    io_s[316] = _zz_io_s_17;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[0:0];
    _zz_io_s_2 <= _zz_io_s[1];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_16 <= _zz_io_s_15[58:0];
    _zz_io_s_17 <= _zz_io_s_15[59];
  end


endmodule

module BADD_541 (
  input      [280:0]  io_a,
  input      [280:0]  io_b,
  input               io_c,
  output reg [281:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [30:0]   _zz__zz_io_s;
  wire       [30:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [59:0]   _zz__zz_io_s_12;
  wire       [59:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [30:0]   _zz_io_s;
  reg        [29:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [59:0]   _zz_io_s_12;
  reg        [58:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[29 : 0]} + {1'b0,io_b[29 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {30'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[93 : 30]} + {1'b0,io_b[93 : 30]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[157 : 94]} + {1'b0,io_b[157 : 94]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[221 : 158]} + {1'b0,io_b[221 : 158]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[280 : 222]} + {1'b0,io_b[280 : 222]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {59'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[29 : 0] = _zz_io_s_1;
    io_s[93 : 30] = _zz_io_s_4;
    io_s[157 : 94] = _zz_io_s_7;
    io_s[221 : 158] = _zz_io_s_10;
    io_s[280 : 222] = _zz_io_s_13;
    io_s[281] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[29:0];
    _zz_io_s_2 <= _zz_io_s[30];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[58:0];
    _zz_io_s_14 <= _zz_io_s_12[59];
  end


endmodule

module BADD_540 (
  input      [276:0]  io_a,
  input      [276:0]  io_b,
  input               io_c,
  output reg [277:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [26:0]   _zz__zz_io_s;
  wire       [26:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [59:0]   _zz__zz_io_s_12;
  wire       [59:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [26:0]   _zz_io_s;
  reg        [25:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [59:0]   _zz_io_s_12;
  reg        [58:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[25 : 0]} + {1'b0,io_b[25 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {26'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[89 : 26]} + {1'b0,io_b[89 : 26]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[153 : 90]} + {1'b0,io_b[153 : 90]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[217 : 154]} + {1'b0,io_b[217 : 154]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[276 : 218]} + {1'b0,io_b[276 : 218]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {59'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[25 : 0] = _zz_io_s_1;
    io_s[89 : 26] = _zz_io_s_4;
    io_s[153 : 90] = _zz_io_s_7;
    io_s[217 : 154] = _zz_io_s_10;
    io_s[276 : 218] = _zz_io_s_13;
    io_s[277] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[25:0];
    _zz_io_s_2 <= _zz_io_s[26];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[58:0];
    _zz_io_s_14 <= _zz_io_s_12[59];
  end


endmodule

module BADD_539 (
  input      [286:0]  io_a,
  input      [286:0]  io_b,
  input               io_c,
  output reg [287:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [36:0]   _zz__zz_io_s;
  wire       [36:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [59:0]   _zz__zz_io_s_12;
  wire       [59:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [36:0]   _zz_io_s;
  reg        [35:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [59:0]   _zz_io_s_12;
  reg        [58:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[35 : 0]} + {1'b0,io_b[35 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {36'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[99 : 36]} + {1'b0,io_b[99 : 36]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[163 : 100]} + {1'b0,io_b[163 : 100]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[227 : 164]} + {1'b0,io_b[227 : 164]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[286 : 228]} + {1'b0,io_b[286 : 228]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {59'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[35 : 0] = _zz_io_s_1;
    io_s[99 : 36] = _zz_io_s_4;
    io_s[163 : 100] = _zz_io_s_7;
    io_s[227 : 164] = _zz_io_s_10;
    io_s[286 : 228] = _zz_io_s_13;
    io_s[287] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[35:0];
    _zz_io_s_2 <= _zz_io_s[36];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[58:0];
    _zz_io_s_14 <= _zz_io_s_12[59];
  end


endmodule

module BADD_538 (
  input      [327:0]  io_a,
  input      [327:0]  io_b,
  input               io_c,
  output reg [328:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [13:0]   _zz__zz_io_s;
  wire       [13:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [59:0]   _zz__zz_io_s_15;
  wire       [59:0]   _zz__zz_io_s_15_1;
  wire       [0:0]    _zz__zz_io_s_15_2;
  wire       [13:0]   _zz_io_s;
  reg        [12:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [59:0]   _zz_io_s_15;
  reg        [58:0]   _zz_io_s_16;
  reg                 _zz_io_s_17;

  assign _zz__zz_io_s = ({1'b0,io_a[12 : 0]} + {1'b0,io_b[12 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {13'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[76 : 13]} + {1'b0,io_b[76 : 13]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[140 : 77]} + {1'b0,io_b[140 : 77]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[204 : 141]} + {1'b0,io_b[204 : 141]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[268 : 205]} + {1'b0,io_b[268 : 205]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[327 : 269]} + {1'b0,io_b[327 : 269]});
  assign _zz__zz_io_s_15_2 = _zz_io_s_14;
  assign _zz__zz_io_s_15_1 = {59'd0, _zz__zz_io_s_15_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[12 : 0] = _zz_io_s_1;
    io_s[76 : 13] = _zz_io_s_4;
    io_s[140 : 77] = _zz_io_s_7;
    io_s[204 : 141] = _zz_io_s_10;
    io_s[268 : 205] = _zz_io_s_13;
    io_s[327 : 269] = _zz_io_s_16;
    io_s[328] = _zz_io_s_17;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[12:0];
    _zz_io_s_2 <= _zz_io_s[13];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_16 <= _zz_io_s_15[58:0];
    _zz_io_s_17 <= _zz_io_s_15[59];
  end


endmodule

module BADD_537 (
  input      [322:0]  io_a,
  input      [322:0]  io_b,
  input               io_c,
  output reg [323:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [8:0]    _zz__zz_io_s;
  wire       [8:0]    _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [59:0]   _zz__zz_io_s_15;
  wire       [59:0]   _zz__zz_io_s_15_1;
  wire       [0:0]    _zz__zz_io_s_15_2;
  wire       [8:0]    _zz_io_s;
  reg        [7:0]    _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [59:0]   _zz_io_s_15;
  reg        [58:0]   _zz_io_s_16;
  reg                 _zz_io_s_17;

  assign _zz__zz_io_s = ({1'b0,io_a[7 : 0]} + {1'b0,io_b[7 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {8'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[71 : 8]} + {1'b0,io_b[71 : 8]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[135 : 72]} + {1'b0,io_b[135 : 72]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[199 : 136]} + {1'b0,io_b[199 : 136]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[263 : 200]} + {1'b0,io_b[263 : 200]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[322 : 264]} + {1'b0,io_b[322 : 264]});
  assign _zz__zz_io_s_15_2 = _zz_io_s_14;
  assign _zz__zz_io_s_15_1 = {59'd0, _zz__zz_io_s_15_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[7 : 0] = _zz_io_s_1;
    io_s[71 : 8] = _zz_io_s_4;
    io_s[135 : 72] = _zz_io_s_7;
    io_s[199 : 136] = _zz_io_s_10;
    io_s[263 : 200] = _zz_io_s_13;
    io_s[322 : 264] = _zz_io_s_16;
    io_s[323] = _zz_io_s_17;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[7:0];
    _zz_io_s_2 <= _zz_io_s[8];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_16 <= _zz_io_s_15[58:0];
    _zz_io_s_17 <= _zz_io_s_15[59];
  end


endmodule

module BADD_536 (
  input      [332:0]  io_a,
  input      [332:0]  io_b,
  input               io_c,
  output reg [333:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [18:0]   _zz__zz_io_s;
  wire       [18:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_3;
  wire       [64:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [64:0]   _zz__zz_io_s_6;
  wire       [64:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [64:0]   _zz__zz_io_s_9;
  wire       [64:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [59:0]   _zz__zz_io_s_15;
  wire       [59:0]   _zz__zz_io_s_15_1;
  wire       [0:0]    _zz__zz_io_s_15_2;
  wire       [18:0]   _zz_io_s;
  reg        [17:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [64:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [64:0]   _zz_io_s_6;
  reg        [63:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [64:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [59:0]   _zz_io_s_15;
  reg        [58:0]   _zz_io_s_16;
  reg                 _zz_io_s_17;

  assign _zz__zz_io_s = ({1'b0,io_a[17 : 0]} + {1'b0,io_b[17 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {18'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[81 : 18]} + {1'b0,io_b[81 : 18]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {64'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[145 : 82]} + {1'b0,io_b[145 : 82]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {64'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[209 : 146]} + {1'b0,io_b[209 : 146]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {64'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[273 : 210]} + {1'b0,io_b[273 : 210]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[332 : 274]} + {1'b0,io_b[332 : 274]});
  assign _zz__zz_io_s_15_2 = _zz_io_s_14;
  assign _zz__zz_io_s_15_1 = {59'd0, _zz__zz_io_s_15_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[17 : 0] = _zz_io_s_1;
    io_s[81 : 18] = _zz_io_s_4;
    io_s[145 : 82] = _zz_io_s_7;
    io_s[209 : 146] = _zz_io_s_10;
    io_s[273 : 210] = _zz_io_s_13;
    io_s[332 : 274] = _zz_io_s_16;
    io_s[333] = _zz_io_s_17;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[17:0];
    _zz_io_s_2 <= _zz_io_s[18];
    _zz_io_s_4 <= _zz_io_s_3[63:0];
    _zz_io_s_5 <= _zz_io_s_3[64];
    _zz_io_s_7 <= _zz_io_s_6[63:0];
    _zz_io_s_8 <= _zz_io_s_6[64];
    _zz_io_s_10 <= _zz_io_s_9[63:0];
    _zz_io_s_11 <= _zz_io_s_9[64];
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_16 <= _zz_io_s_15[58:0];
    _zz_io_s_17 <= _zz_io_s_15[59];
  end


endmodule

module BADD_535 (
  input      [189:0]  io_a,
  input      [189:0]  io_b,
  input               io_c,
  output reg [190:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [189:0]  _zz__zz_io_s_1;
  wire       [64:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [189:0]  _zz__zz_io_s_4;
  wire       [64:0]   _zz__zz_io_s_5;
  wire       [64:0]   _zz__zz_io_s_5_1;
  wire       [0:0]    _zz__zz_io_s_5_2;
  wire       [189:0]  _zz__zz_io_s_10;
  wire       [62:0]   _zz__zz_io_s_12;
  wire       [62:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  wire       [64:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [61:0]   _zz_io_s_8;
  reg        [61:0]   _zz_io_s_9;
  reg        [61:0]   _zz_io_s_10;
  reg        [61:0]   _zz_io_s_11;
  wire       [62:0]   _zz_io_s_12;
  reg        [61:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,_zz__zz_io_s_1[63 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {64'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_4 = (~ io_b);
  assign _zz__zz_io_s_5 = ({1'b0,_zz_io_s_3} + {1'b0,_zz_io_s_4});
  assign _zz__zz_io_s_5_2 = _zz_io_s_2;
  assign _zz__zz_io_s_5_1 = {64'd0, _zz__zz_io_s_5_2};
  assign _zz__zz_io_s_10 = (~ io_b);
  assign _zz__zz_io_s_12 = ({1'b0,_zz_io_s_9} + {1'b0,_zz_io_s_11});
  assign _zz__zz_io_s_12_2 = _zz_io_s_7;
  assign _zz__zz_io_s_12_1 = {62'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_1;
    io_s[127 : 64] = _zz_io_s_6;
    io_s[189 : 128] = _zz_io_s_13;
    io_s[190] = (! _zz_io_s_14);
  end

  assign _zz_io_s_5 = (_zz__zz_io_s_5 + _zz__zz_io_s_5_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s[64];
    _zz_io_s_3 <= io_a[127 : 64];
    _zz_io_s_4 <= _zz__zz_io_s_4[127 : 64];
    _zz_io_s_6 <= _zz_io_s_5[63:0];
    _zz_io_s_7 <= _zz_io_s_5[64];
    _zz_io_s_8 <= io_a[189 : 128];
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= _zz__zz_io_s_10[189 : 128];
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_13 <= _zz_io_s_12[61:0];
    _zz_io_s_14 <= _zz_io_s_12[62];
  end


endmodule

module BADD_534 (
  input      [272:0]  io_a,
  input      [272:0]  io_b,
  input               io_c,
  output reg [273:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [64:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_5;
  wire       [64:0]   _zz__zz_io_s_5_1;
  wire       [0:0]    _zz__zz_io_s_5_2;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [17:0]   _zz__zz_io_s_32;
  wire       [17:0]   _zz__zz_io_s_32_1;
  wire       [0:0]    _zz__zz_io_s_32_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  wire       [64:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  reg        [16:0]   _zz_io_s_24;
  reg        [16:0]   _zz_io_s_25;
  reg        [16:0]   _zz_io_s_26;
  reg        [16:0]   _zz_io_s_27;
  reg        [16:0]   _zz_io_s_28;
  reg        [16:0]   _zz_io_s_29;
  reg        [16:0]   _zz_io_s_30;
  reg        [16:0]   _zz_io_s_31;
  wire       [17:0]   _zz_io_s_32;
  reg        [16:0]   _zz_io_s_33;
  reg                 _zz_io_s_34;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,io_b[63 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {64'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_5 = ({1'b0,_zz_io_s_3} + {1'b0,_zz_io_s_4});
  assign _zz__zz_io_s_5_2 = _zz_io_s_2;
  assign _zz__zz_io_s_5_1 = {64'd0, _zz__zz_io_s_5_2};
  assign _zz__zz_io_s_12 = ({1'b0,_zz_io_s_9} + {1'b0,_zz_io_s_11});
  assign _zz__zz_io_s_12_2 = _zz_io_s_7;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_17} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_14;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_32 = ({1'b0,_zz_io_s_27} + {1'b0,_zz_io_s_31});
  assign _zz__zz_io_s_32_2 = _zz_io_s_23;
  assign _zz__zz_io_s_32_1 = {17'd0, _zz__zz_io_s_32_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_1;
    io_s[127 : 64] = _zz_io_s_6;
    io_s[191 : 128] = _zz_io_s_13;
    io_s[255 : 192] = _zz_io_s_22;
    io_s[272 : 256] = _zz_io_s_33;
    io_s[273] = _zz_io_s_34;
  end

  assign _zz_io_s_5 = (_zz__zz_io_s_5 + _zz__zz_io_s_5_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_32 = (_zz__zz_io_s_32 + _zz__zz_io_s_32_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s[64];
    _zz_io_s_3 <= io_a[127 : 64];
    _zz_io_s_4 <= io_b[127 : 64];
    _zz_io_s_6 <= _zz_io_s_5[63:0];
    _zz_io_s_7 <= _zz_io_s_5[64];
    _zz_io_s_8 <= io_a[191 : 128];
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= io_b[191 : 128];
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_15 <= io_a[255 : 192];
    _zz_io_s_16 <= _zz_io_s_15;
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= io_b[255 : 192];
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_21[64];
    _zz_io_s_24 <= io_a[272 : 256];
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_25;
    _zz_io_s_27 <= _zz_io_s_26;
    _zz_io_s_28 <= io_b[272 : 256];
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz_io_s_29;
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_33 <= _zz_io_s_32[16:0];
    _zz_io_s_34 <= _zz_io_s_32[17];
  end


endmodule

module BADD_533 (
  input      [332:0]  io_a,
  input      [332:0]  io_b,
  input               io_c,
  output reg [333:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [64:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_5;
  wire       [64:0]   _zz__zz_io_s_5_1;
  wire       [0:0]    _zz__zz_io_s_5_2;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [64:0]   _zz__zz_io_s_32;
  wire       [64:0]   _zz__zz_io_s_32_1;
  wire       [0:0]    _zz__zz_io_s_32_2;
  wire       [13:0]   _zz__zz_io_s_45;
  wire       [13:0]   _zz__zz_io_s_45_1;
  wire       [0:0]    _zz__zz_io_s_45_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  wire       [64:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg        [63:0]   _zz_io_s_25;
  reg        [63:0]   _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg        [63:0]   _zz_io_s_29;
  reg        [63:0]   _zz_io_s_30;
  reg        [63:0]   _zz_io_s_31;
  wire       [64:0]   _zz_io_s_32;
  reg        [63:0]   _zz_io_s_33;
  reg                 _zz_io_s_34;
  reg        [12:0]   _zz_io_s_35;
  reg        [12:0]   _zz_io_s_36;
  reg        [12:0]   _zz_io_s_37;
  reg        [12:0]   _zz_io_s_38;
  reg        [12:0]   _zz_io_s_39;
  reg        [12:0]   _zz_io_s_40;
  reg        [12:0]   _zz_io_s_41;
  reg        [12:0]   _zz_io_s_42;
  reg        [12:0]   _zz_io_s_43;
  reg        [12:0]   _zz_io_s_44;
  wire       [13:0]   _zz_io_s_45;
  reg        [12:0]   _zz_io_s_46;
  reg                 _zz_io_s_47;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,io_b[63 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {64'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_5 = ({1'b0,_zz_io_s_3} + {1'b0,_zz_io_s_4});
  assign _zz__zz_io_s_5_2 = _zz_io_s_2;
  assign _zz__zz_io_s_5_1 = {64'd0, _zz__zz_io_s_5_2};
  assign _zz__zz_io_s_12 = ({1'b0,_zz_io_s_9} + {1'b0,_zz_io_s_11});
  assign _zz__zz_io_s_12_2 = _zz_io_s_7;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_17} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_14;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_32 = ({1'b0,_zz_io_s_27} + {1'b0,_zz_io_s_31});
  assign _zz__zz_io_s_32_2 = _zz_io_s_23;
  assign _zz__zz_io_s_32_1 = {64'd0, _zz__zz_io_s_32_2};
  assign _zz__zz_io_s_45 = ({1'b0,_zz_io_s_39} + {1'b0,_zz_io_s_44});
  assign _zz__zz_io_s_45_2 = _zz_io_s_34;
  assign _zz__zz_io_s_45_1 = {13'd0, _zz__zz_io_s_45_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_1;
    io_s[127 : 64] = _zz_io_s_6;
    io_s[191 : 128] = _zz_io_s_13;
    io_s[255 : 192] = _zz_io_s_22;
    io_s[319 : 256] = _zz_io_s_33;
    io_s[332 : 320] = _zz_io_s_46;
    io_s[333] = _zz_io_s_47;
  end

  assign _zz_io_s_5 = (_zz__zz_io_s_5 + _zz__zz_io_s_5_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_32 = (_zz__zz_io_s_32 + _zz__zz_io_s_32_1);
  assign _zz_io_s_45 = (_zz__zz_io_s_45 + _zz__zz_io_s_45_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s[64];
    _zz_io_s_3 <= io_a[127 : 64];
    _zz_io_s_4 <= io_b[127 : 64];
    _zz_io_s_6 <= _zz_io_s_5[63:0];
    _zz_io_s_7 <= _zz_io_s_5[64];
    _zz_io_s_8 <= io_a[191 : 128];
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= io_b[191 : 128];
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_15 <= io_a[255 : 192];
    _zz_io_s_16 <= _zz_io_s_15;
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= io_b[255 : 192];
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_21[64];
    _zz_io_s_24 <= io_a[319 : 256];
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_25;
    _zz_io_s_27 <= _zz_io_s_26;
    _zz_io_s_28 <= io_b[319 : 256];
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz_io_s_29;
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_33 <= _zz_io_s_32[63:0];
    _zz_io_s_34 <= _zz_io_s_32[64];
    _zz_io_s_35 <= io_a[332 : 320];
    _zz_io_s_36 <= _zz_io_s_35;
    _zz_io_s_37 <= _zz_io_s_36;
    _zz_io_s_38 <= _zz_io_s_37;
    _zz_io_s_39 <= _zz_io_s_38;
    _zz_io_s_40 <= io_b[332 : 320];
    _zz_io_s_41 <= _zz_io_s_40;
    _zz_io_s_42 <= _zz_io_s_41;
    _zz_io_s_43 <= _zz_io_s_42;
    _zz_io_s_44 <= _zz_io_s_43;
    _zz_io_s_46 <= _zz_io_s_45[12:0];
    _zz_io_s_47 <= _zz_io_s_45[13];
  end


endmodule

module BADD_532 (
  input      [322:0]  io_a,
  input      [322:0]  io_b,
  input               io_c,
  output reg [323:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [64:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_5;
  wire       [64:0]   _zz__zz_io_s_5_1;
  wire       [0:0]    _zz__zz_io_s_5_2;
  wire       [64:0]   _zz__zz_io_s_12;
  wire       [64:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [64:0]   _zz__zz_io_s_32;
  wire       [64:0]   _zz__zz_io_s_32_1;
  wire       [0:0]    _zz__zz_io_s_32_2;
  wire       [3:0]    _zz__zz_io_s_45;
  wire       [3:0]    _zz__zz_io_s_45_1;
  wire       [0:0]    _zz__zz_io_s_45_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  wire       [64:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  reg        [63:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  wire       [64:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  reg        [63:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg        [63:0]   _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg        [63:0]   _zz_io_s_25;
  reg        [63:0]   _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg        [63:0]   _zz_io_s_29;
  reg        [63:0]   _zz_io_s_30;
  reg        [63:0]   _zz_io_s_31;
  wire       [64:0]   _zz_io_s_32;
  reg        [63:0]   _zz_io_s_33;
  reg                 _zz_io_s_34;
  reg        [2:0]    _zz_io_s_35;
  reg        [2:0]    _zz_io_s_36;
  reg        [2:0]    _zz_io_s_37;
  reg        [2:0]    _zz_io_s_38;
  reg        [2:0]    _zz_io_s_39;
  reg        [2:0]    _zz_io_s_40;
  reg        [2:0]    _zz_io_s_41;
  reg        [2:0]    _zz_io_s_42;
  reg        [2:0]    _zz_io_s_43;
  reg        [2:0]    _zz_io_s_44;
  wire       [3:0]    _zz_io_s_45;
  reg        [2:0]    _zz_io_s_46;
  reg                 _zz_io_s_47;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,io_b[63 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {64'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_5 = ({1'b0,_zz_io_s_3} + {1'b0,_zz_io_s_4});
  assign _zz__zz_io_s_5_2 = _zz_io_s_2;
  assign _zz__zz_io_s_5_1 = {64'd0, _zz__zz_io_s_5_2};
  assign _zz__zz_io_s_12 = ({1'b0,_zz_io_s_9} + {1'b0,_zz_io_s_11});
  assign _zz__zz_io_s_12_2 = _zz_io_s_7;
  assign _zz__zz_io_s_12_1 = {64'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_21 = ({1'b0,_zz_io_s_17} + {1'b0,_zz_io_s_20});
  assign _zz__zz_io_s_21_2 = _zz_io_s_14;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_32 = ({1'b0,_zz_io_s_27} + {1'b0,_zz_io_s_31});
  assign _zz__zz_io_s_32_2 = _zz_io_s_23;
  assign _zz__zz_io_s_32_1 = {64'd0, _zz__zz_io_s_32_2};
  assign _zz__zz_io_s_45 = ({1'b0,_zz_io_s_39} + {1'b0,_zz_io_s_44});
  assign _zz__zz_io_s_45_2 = _zz_io_s_34;
  assign _zz__zz_io_s_45_1 = {3'd0, _zz__zz_io_s_45_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_1;
    io_s[127 : 64] = _zz_io_s_6;
    io_s[191 : 128] = _zz_io_s_13;
    io_s[255 : 192] = _zz_io_s_22;
    io_s[319 : 256] = _zz_io_s_33;
    io_s[322 : 320] = _zz_io_s_46;
    io_s[323] = _zz_io_s_47;
  end

  assign _zz_io_s_5 = (_zz__zz_io_s_5 + _zz__zz_io_s_5_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_32 = (_zz__zz_io_s_32 + _zz__zz_io_s_32_1);
  assign _zz_io_s_45 = (_zz__zz_io_s_45 + _zz__zz_io_s_45_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s[64];
    _zz_io_s_3 <= io_a[127 : 64];
    _zz_io_s_4 <= io_b[127 : 64];
    _zz_io_s_6 <= _zz_io_s_5[63:0];
    _zz_io_s_7 <= _zz_io_s_5[64];
    _zz_io_s_8 <= io_a[191 : 128];
    _zz_io_s_9 <= _zz_io_s_8;
    _zz_io_s_10 <= io_b[191 : 128];
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_13 <= _zz_io_s_12[63:0];
    _zz_io_s_14 <= _zz_io_s_12[64];
    _zz_io_s_15 <= io_a[255 : 192];
    _zz_io_s_16 <= _zz_io_s_15;
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= io_b[255 : 192];
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_19;
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_21[64];
    _zz_io_s_24 <= io_a[319 : 256];
    _zz_io_s_25 <= _zz_io_s_24;
    _zz_io_s_26 <= _zz_io_s_25;
    _zz_io_s_27 <= _zz_io_s_26;
    _zz_io_s_28 <= io_b[319 : 256];
    _zz_io_s_29 <= _zz_io_s_28;
    _zz_io_s_30 <= _zz_io_s_29;
    _zz_io_s_31 <= _zz_io_s_30;
    _zz_io_s_33 <= _zz_io_s_32[63:0];
    _zz_io_s_34 <= _zz_io_s_32[64];
    _zz_io_s_35 <= io_a[322 : 320];
    _zz_io_s_36 <= _zz_io_s_35;
    _zz_io_s_37 <= _zz_io_s_36;
    _zz_io_s_38 <= _zz_io_s_37;
    _zz_io_s_39 <= _zz_io_s_38;
    _zz_io_s_40 <= io_b[322 : 320];
    _zz_io_s_41 <= _zz_io_s_40;
    _zz_io_s_42 <= _zz_io_s_41;
    _zz_io_s_43 <= _zz_io_s_42;
    _zz_io_s_44 <= _zz_io_s_43;
    _zz_io_s_46 <= _zz_io_s_45[2:0];
    _zz_io_s_47 <= _zz_io_s_45[3];
  end


endmodule

//KaratsubaCore_16 replaced by KaratsubaCore_17

module KaratsubaCore_17 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_a_2,
  input      [47:0]   io_a_3,
  input      [47:0]   io_a_4,
  input      [47:0]   io_a_5,
  input      [47:0]   io_a_6,
  input      [47:0]   io_a_7,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  input      [47:0]   io_b_2,
  input      [47:0]   io_b_3,
  input      [47:0]   io_b_4,
  input      [47:0]   io_b_5,
  input      [47:0]   io_b_6,
  input      [47:0]   io_b_7,
  output reg [767:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [384:0]  karatsuba_add2_io_a;
  wire       [575:0]  karatsuba_noExtend_add3_io_a;
  reg        [575:0]  karatsuba_noExtend_add3_io_b;
  wire       [383:0]  karatsuba_lsbMul_io_p;
  wire       [385:0]  karatsuba_midMul_io_p;
  wire       [383:0]  karatsuba_msbMul_io_p;
  wire       [384:0]  karatsuba_add1_io_s;
  wire       [385:0]  karatsuba_add2_io_s;
  wire       [576:0]  karatsuba_noExtend_add3_io_s;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_a_1;
  reg        [48:0]   _zz_io_a_2;
  reg        [48:0]   _zz_io_a_3;
  reg        [48:0]   _zz_io_b_0;
  reg        [48:0]   _zz_io_b_1;
  reg        [48:0]   _zz_io_b_2;
  reg        [48:0]   _zz_io_b_3;
  reg        [384:0]  core_karatsuba_add1_io_s_delay_1;
  reg        [384:0]  _zz_io_a;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_1;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_2;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_3;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_4;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_5;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_6;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_7;
  reg        [383:0]  core_karatsuba_msbMul_io_p_delay_8;
  reg        [191:0]  _zz_io_p;

  KaratsubaCore_69 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]                ), //i
    .io_a_1 (io_a_1[47:0]                ), //i
    .io_a_2 (io_a_2[47:0]                ), //i
    .io_a_3 (io_a_3[47:0]                ), //i
    .io_b_0 (io_b_0[47:0]                ), //i
    .io_b_1 (io_b_1[47:0]                ), //i
    .io_b_2 (io_b_2[47:0]                ), //i
    .io_b_3 (io_b_3[47:0]                ), //i
    .io_p   (karatsuba_lsbMul_io_p[383:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_70 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]            ), //i
    .io_a_1 (_zz_io_a_1[48:0]            ), //i
    .io_a_2 (_zz_io_a_2[48:0]            ), //i
    .io_a_3 (_zz_io_a_3[48:0]            ), //i
    .io_b_0 (_zz_io_b_0[48:0]            ), //i
    .io_b_1 (_zz_io_b_1[48:0]            ), //i
    .io_b_2 (_zz_io_b_2[48:0]            ), //i
    .io_b_3 (_zz_io_b_3[48:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[385:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_71 karatsuba_msbMul (
    .io_a_0 (io_a_4[47:0]                ), //i
    .io_a_1 (io_a_5[47:0]                ), //i
    .io_a_2 (io_a_6[47:0]                ), //i
    .io_a_3 (io_a_7[47:0]                ), //i
    .io_b_0 (io_b_4[47:0]                ), //i
    .io_b_1 (io_b_5[47:0]                ), //i
    .io_b_2 (io_b_6[47:0]                ), //i
    .io_b_3 (io_b_7[47:0]                ), //i
    .io_p   (karatsuba_msbMul_io_p[383:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_654 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[383:0]), //i
    .io_b   (karatsuba_msbMul_io_p[383:0]), //i
    .io_c   (1'b0                        ), //i
    .io_s   (karatsuba_add1_io_s[384:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_655 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[384:0]             ), //i
    .io_b   (core_karatsuba_add1_io_s_delay_1[384:0]), //i
    .io_c   (1'b1                                   ), //i
    .io_s   (karatsuba_add2_io_s[385:0]             ), //o
    .clk    (clk                                    ), //i
    .resetn (resetn                                 )  //i
  );
  BADD_656 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[575:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[575:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[576:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[384:0];
  assign karatsuba_noExtend_add3_io_a = {191'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[191 : 0] = (karatsuba_lsbMul_io_p >>> 192);
    karatsuba_noExtend_add3_io_b[575 : 192] = core_karatsuba_msbMul_io_p_delay_8;
  end

  always @(*) begin
    io_p[191 : 0] = _zz_io_p;
    io_p[767 : 192] = karatsuba_noExtend_add3_io_s[575:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_4});
    _zz_io_a_1 <= ({1'b0,io_a_1} + {1'b0,io_a_5});
    _zz_io_a_2 <= ({1'b0,io_a_2} + {1'b0,io_a_6});
    _zz_io_a_3 <= ({1'b0,io_a_3} + {1'b0,io_a_7});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_4});
    _zz_io_b_1 <= ({1'b0,io_b_1} + {1'b0,io_b_5});
    _zz_io_b_2 <= ({1'b0,io_b_2} + {1'b0,io_b_6});
    _zz_io_b_3 <= ({1'b0,io_b_3} + {1'b0,io_b_7});
    core_karatsuba_add1_io_s_delay_1 <= karatsuba_add1_io_s;
    _zz_io_a <= karatsuba_add2_io_s[384:0];
    core_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    core_karatsuba_msbMul_io_p_delay_2 <= core_karatsuba_msbMul_io_p_delay_1;
    core_karatsuba_msbMul_io_p_delay_3 <= core_karatsuba_msbMul_io_p_delay_2;
    core_karatsuba_msbMul_io_p_delay_4 <= core_karatsuba_msbMul_io_p_delay_3;
    core_karatsuba_msbMul_io_p_delay_5 <= core_karatsuba_msbMul_io_p_delay_4;
    core_karatsuba_msbMul_io_p_delay_6 <= core_karatsuba_msbMul_io_p_delay_5;
    core_karatsuba_msbMul_io_p_delay_7 <= core_karatsuba_msbMul_io_p_delay_6;
    core_karatsuba_msbMul_io_p_delay_8 <= core_karatsuba_msbMul_io_p_delay_7;
    _zz_io_p <= karatsuba_lsbMul_io_p[191 : 0];
  end


endmodule

//BADD_594 replaced by BADD_650

//BADD_597 replaced by BADD_656

//BADD_596 replaced by BADD_655

//BADD_595 replaced by BADD_654

//KaratsubaCore_20 replaced by KaratsubaCore_71

//KaratsubaCore_19 replaced by KaratsubaCore_70

//KaratsubaCore_18 replaced by KaratsubaCore_69

//BADD_600 replaced by BADD_656

//BADD_599 replaced by BADD_655

//BADD_598 replaced by BADD_654

//KaratsubaCore_23 replaced by KaratsubaCore_71

//KaratsubaCore_22 replaced by KaratsubaCore_70

//KaratsubaCore_21 replaced by KaratsubaCore_69

//BADD_601 replaced by BADD_650

//BADD_604 replaced by BADD_656

//BADD_603 replaced by BADD_655

//BADD_602 replaced by BADD_654

//KaratsubaCore_26 replaced by KaratsubaCore_71

//KaratsubaCore_25 replaced by KaratsubaCore_70

//KaratsubaCore_24 replaced by KaratsubaCore_69

//BADD_607 replaced by BADD_656

//BADD_606 replaced by BADD_655

//BADD_605 replaced by BADD_654

//KaratsubaCore_29 replaced by KaratsubaCore_71

//KaratsubaCore_28 replaced by KaratsubaCore_70

//KaratsubaCore_27 replaced by KaratsubaCore_69

//BADD_608 replaced by BADD_650

//BADD_611 replaced by BADD_656

//BADD_610 replaced by BADD_655

//BADD_609 replaced by BADD_654

//KaratsubaCore_32 replaced by KaratsubaCore_71

//KaratsubaCore_31 replaced by KaratsubaCore_70

//KaratsubaCore_30 replaced by KaratsubaCore_69

//BADD_614 replaced by BADD_656

//BADD_613 replaced by BADD_655

//BADD_612 replaced by BADD_654

//KaratsubaCore_35 replaced by KaratsubaCore_71

//KaratsubaCore_34 replaced by KaratsubaCore_70

//KaratsubaCore_33 replaced by KaratsubaCore_69

//BADD_615 replaced by BADD_650

//BADD_618 replaced by BADD_656

//BADD_617 replaced by BADD_655

//BADD_616 replaced by BADD_654

//KaratsubaCore_38 replaced by KaratsubaCore_71

//KaratsubaCore_37 replaced by KaratsubaCore_70

//KaratsubaCore_36 replaced by KaratsubaCore_69

//BADD_621 replaced by BADD_656

//BADD_620 replaced by BADD_655

//BADD_619 replaced by BADD_654

//KaratsubaCore_41 replaced by KaratsubaCore_71

//KaratsubaCore_40 replaced by KaratsubaCore_70

//KaratsubaCore_39 replaced by KaratsubaCore_69

//BADD_622 replaced by BADD_650

//BADD_625 replaced by BADD_656

//BADD_624 replaced by BADD_655

//BADD_623 replaced by BADD_654

//KaratsubaCore_44 replaced by KaratsubaCore_71

//KaratsubaCore_43 replaced by KaratsubaCore_70

//KaratsubaCore_42 replaced by KaratsubaCore_69

//BADD_628 replaced by BADD_656

//BADD_627 replaced by BADD_655

//BADD_626 replaced by BADD_654

//KaratsubaCore_47 replaced by KaratsubaCore_71

//KaratsubaCore_46 replaced by KaratsubaCore_70

//KaratsubaCore_45 replaced by KaratsubaCore_69

//BADD_629 replaced by BADD_650

//BADD_632 replaced by BADD_656

//BADD_631 replaced by BADD_655

//BADD_630 replaced by BADD_654

//KaratsubaCore_50 replaced by KaratsubaCore_71

//KaratsubaCore_49 replaced by KaratsubaCore_70

//KaratsubaCore_48 replaced by KaratsubaCore_69

//BADD_635 replaced by BADD_656

//BADD_634 replaced by BADD_655

//BADD_633 replaced by BADD_654

//KaratsubaCore_53 replaced by KaratsubaCore_71

//KaratsubaCore_52 replaced by KaratsubaCore_70

//KaratsubaCore_51 replaced by KaratsubaCore_69

//BADD_636 replaced by BADD_650

//BADD_639 replaced by BADD_656

//BADD_638 replaced by BADD_655

//BADD_637 replaced by BADD_654

//KaratsubaCore_56 replaced by KaratsubaCore_71

//KaratsubaCore_55 replaced by KaratsubaCore_70

//KaratsubaCore_54 replaced by KaratsubaCore_69

//BADD_642 replaced by BADD_656

//BADD_641 replaced by BADD_655

//BADD_640 replaced by BADD_654

//KaratsubaCore_59 replaced by KaratsubaCore_71

//KaratsubaCore_58 replaced by KaratsubaCore_70

//KaratsubaCore_57 replaced by KaratsubaCore_69

//BADD_643 replaced by BADD_650

//BADD_646 replaced by BADD_656

//BADD_645 replaced by BADD_655

//BADD_644 replaced by BADD_654

//KaratsubaCore_62 replaced by KaratsubaCore_71

//KaratsubaCore_61 replaced by KaratsubaCore_70

//KaratsubaCore_60 replaced by KaratsubaCore_69

//BADD_649 replaced by BADD_656

//BADD_648 replaced by BADD_655

//BADD_647 replaced by BADD_654

//KaratsubaCore_65 replaced by KaratsubaCore_71

//KaratsubaCore_64 replaced by KaratsubaCore_70

//KaratsubaCore_63 replaced by KaratsubaCore_69

module BADD_650 (
  input      [377:0]  io_a,
  input      [377:0]  io_b,
  input               io_c,
  output reg [378:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [64:0]   _zz__zz_io_s;
  wire       [64:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [64:0]   _zz__zz_io_s_8;
  wire       [64:0]   _zz__zz_io_s_8_1;
  wire       [0:0]    _zz__zz_io_s_8_2;
  wire       [64:0]   _zz__zz_io_s_15;
  wire       [64:0]   _zz__zz_io_s_15_1;
  wire       [0:0]    _zz__zz_io_s_15_2;
  wire       [64:0]   _zz__zz_io_s_21;
  wire       [64:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [64:0]   _zz__zz_io_s_26;
  wire       [64:0]   _zz__zz_io_s_26_1;
  wire       [0:0]    _zz__zz_io_s_26_2;
  wire       [58:0]   _zz__zz_io_s_30;
  wire       [58:0]   _zz__zz_io_s_30_1;
  wire       [0:0]    _zz__zz_io_s_30_2;
  wire       [64:0]   _zz_io_s;
  reg        [63:0]   _zz_io_s_1;
  reg        [63:0]   _zz_io_s_2;
  reg        [63:0]   _zz_io_s_3;
  reg        [63:0]   _zz_io_s_4;
  reg        [63:0]   _zz_io_s_5;
  reg        [63:0]   _zz_io_s_6;
  reg                 _zz_io_s_7;
  wire       [64:0]   _zz_io_s_8;
  reg        [63:0]   _zz_io_s_9;
  reg        [63:0]   _zz_io_s_10;
  reg        [63:0]   _zz_io_s_11;
  reg        [63:0]   _zz_io_s_12;
  reg        [63:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [64:0]   _zz_io_s_15;
  reg        [63:0]   _zz_io_s_16;
  reg        [63:0]   _zz_io_s_17;
  reg        [63:0]   _zz_io_s_18;
  reg        [63:0]   _zz_io_s_19;
  reg                 _zz_io_s_20;
  wire       [64:0]   _zz_io_s_21;
  reg        [63:0]   _zz_io_s_22;
  reg        [63:0]   _zz_io_s_23;
  reg        [63:0]   _zz_io_s_24;
  reg                 _zz_io_s_25;
  wire       [64:0]   _zz_io_s_26;
  reg        [63:0]   _zz_io_s_27;
  reg        [63:0]   _zz_io_s_28;
  reg                 _zz_io_s_29;
  wire       [58:0]   _zz_io_s_30;
  reg        [57:0]   _zz_io_s_31;
  reg                 _zz_io_s_32;

  assign _zz__zz_io_s = ({1'b0,io_a[63 : 0]} + {1'b0,io_b[63 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {64'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_8 = ({1'b0,io_a[127 : 64]} + {1'b0,io_b[127 : 64]});
  assign _zz__zz_io_s_8_2 = _zz_io_s_7;
  assign _zz__zz_io_s_8_1 = {64'd0, _zz__zz_io_s_8_2};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[191 : 128]} + {1'b0,io_b[191 : 128]});
  assign _zz__zz_io_s_15_2 = _zz_io_s_14;
  assign _zz__zz_io_s_15_1 = {64'd0, _zz__zz_io_s_15_2};
  assign _zz__zz_io_s_21 = ({1'b0,io_a[255 : 192]} + {1'b0,io_b[255 : 192]});
  assign _zz__zz_io_s_21_2 = _zz_io_s_20;
  assign _zz__zz_io_s_21_1 = {64'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_26 = ({1'b0,io_a[319 : 256]} + {1'b0,io_b[319 : 256]});
  assign _zz__zz_io_s_26_2 = _zz_io_s_25;
  assign _zz__zz_io_s_26_1 = {64'd0, _zz__zz_io_s_26_2};
  assign _zz__zz_io_s_30 = ({1'b0,io_a[377 : 320]} + {1'b0,io_b[377 : 320]});
  assign _zz__zz_io_s_30_2 = _zz_io_s_29;
  assign _zz__zz_io_s_30_1 = {58'd0, _zz__zz_io_s_30_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[63 : 0] = _zz_io_s_6;
    io_s[127 : 64] = _zz_io_s_13;
    io_s[191 : 128] = _zz_io_s_19;
    io_s[255 : 192] = _zz_io_s_24;
    io_s[319 : 256] = _zz_io_s_28;
    io_s[377 : 320] = _zz_io_s_31;
    io_s[378] = _zz_io_s_32;
  end

  assign _zz_io_s_8 = (_zz__zz_io_s_8 + _zz__zz_io_s_8_1);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_26 = (_zz__zz_io_s_26 + _zz__zz_io_s_26_1);
  assign _zz_io_s_30 = (_zz__zz_io_s_30 + _zz__zz_io_s_30_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[63:0];
    _zz_io_s_2 <= _zz_io_s_1;
    _zz_io_s_3 <= _zz_io_s_2;
    _zz_io_s_4 <= _zz_io_s_3;
    _zz_io_s_5 <= _zz_io_s_4;
    _zz_io_s_6 <= _zz_io_s_5;
    _zz_io_s_7 <= _zz_io_s[64];
    _zz_io_s_9 <= _zz_io_s_8[63:0];
    _zz_io_s_10 <= _zz_io_s_9;
    _zz_io_s_11 <= _zz_io_s_10;
    _zz_io_s_12 <= _zz_io_s_11;
    _zz_io_s_13 <= _zz_io_s_12;
    _zz_io_s_14 <= _zz_io_s_8[64];
    _zz_io_s_16 <= _zz_io_s_15[63:0];
    _zz_io_s_17 <= _zz_io_s_16;
    _zz_io_s_18 <= _zz_io_s_17;
    _zz_io_s_19 <= _zz_io_s_18;
    _zz_io_s_20 <= _zz_io_s_15[64];
    _zz_io_s_22 <= _zz_io_s_21[63:0];
    _zz_io_s_23 <= _zz_io_s_22;
    _zz_io_s_24 <= _zz_io_s_23;
    _zz_io_s_25 <= _zz_io_s_21[64];
    _zz_io_s_27 <= _zz_io_s_26[63:0];
    _zz_io_s_28 <= _zz_io_s_27;
    _zz_io_s_29 <= _zz_io_s_26[64];
    _zz_io_s_31 <= _zz_io_s_30[57:0];
    _zz_io_s_32 <= _zz_io_s_30[58];
  end


endmodule

//BADD_653 replaced by BADD_656

//BADD_652 replaced by BADD_655

//BADD_651 replaced by BADD_654

//KaratsubaCore_68 replaced by KaratsubaCore_71

//KaratsubaCore_67 replaced by KaratsubaCore_70

//KaratsubaCore_66 replaced by KaratsubaCore_69

module BADD_656 (
  input      [575:0]  io_a,
  input      [575:0]  io_b,
  input               io_c,
  output reg [576:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [48:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [48:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [48:0]   _zz__zz_io_s_12;
  wire       [48:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [48:0]   _zz__zz_io_s_15;
  wire       [48:0]   _zz__zz_io_s_15_1;
  wire       [0:0]    _zz__zz_io_s_15_2;
  wire       [48:0]   _zz__zz_io_s_18;
  wire       [48:0]   _zz__zz_io_s_18_1;
  wire       [0:0]    _zz__zz_io_s_18_2;
  wire       [48:0]   _zz__zz_io_s_21;
  wire       [48:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [48:0]   _zz__zz_io_s_24;
  wire       [48:0]   _zz__zz_io_s_24_1;
  wire       [0:0]    _zz__zz_io_s_24_2;
  wire       [48:0]   _zz__zz_io_s_27;
  wire       [48:0]   _zz__zz_io_s_27_1;
  wire       [0:0]    _zz__zz_io_s_27_2;
  wire       [48:0]   _zz__zz_io_s_30;
  wire       [48:0]   _zz__zz_io_s_30_1;
  wire       [0:0]    _zz__zz_io_s_30_2;
  wire       [48:0]   _zz__zz_io_s_33;
  wire       [48:0]   _zz__zz_io_s_33_1;
  wire       [0:0]    _zz__zz_io_s_33_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [48:0]   _zz_io_s_12;
  reg        [47:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [48:0]   _zz_io_s_15;
  reg        [47:0]   _zz_io_s_16;
  reg                 _zz_io_s_17;
  wire       [48:0]   _zz_io_s_18;
  reg        [47:0]   _zz_io_s_19;
  reg                 _zz_io_s_20;
  wire       [48:0]   _zz_io_s_21;
  reg        [47:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  wire       [48:0]   _zz_io_s_24;
  reg        [47:0]   _zz_io_s_25;
  reg                 _zz_io_s_26;
  wire       [48:0]   _zz_io_s_27;
  reg        [47:0]   _zz_io_s_28;
  reg                 _zz_io_s_29;
  wire       [48:0]   _zz_io_s_30;
  reg        [47:0]   _zz_io_s_31;
  reg                 _zz_io_s_32;
  wire       [48:0]   _zz_io_s_33;
  reg        [47:0]   _zz_io_s_34;
  reg                 _zz_io_s_35;
  reg                 _zz_io_s_36;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,io_b[143 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {48'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,io_b[191 : 144]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {48'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[239 : 192]} + {1'b0,io_b[239 : 192]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {48'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[287 : 240]} + {1'b0,io_b[287 : 240]});
  assign _zz__zz_io_s_15_2 = _zz_io_s_14;
  assign _zz__zz_io_s_15_1 = {48'd0, _zz__zz_io_s_15_2};
  assign _zz__zz_io_s_18 = ({1'b0,io_a[335 : 288]} + {1'b0,io_b[335 : 288]});
  assign _zz__zz_io_s_18_2 = _zz_io_s_17;
  assign _zz__zz_io_s_18_1 = {48'd0, _zz__zz_io_s_18_2};
  assign _zz__zz_io_s_21 = ({1'b0,io_a[383 : 336]} + {1'b0,io_b[383 : 336]});
  assign _zz__zz_io_s_21_2 = _zz_io_s_20;
  assign _zz__zz_io_s_21_1 = {48'd0, _zz__zz_io_s_21_2};
  assign _zz__zz_io_s_24 = ({1'b0,io_a[431 : 384]} + {1'b0,io_b[431 : 384]});
  assign _zz__zz_io_s_24_2 = _zz_io_s_23;
  assign _zz__zz_io_s_24_1 = {48'd0, _zz__zz_io_s_24_2};
  assign _zz__zz_io_s_27 = ({1'b0,io_a[479 : 432]} + {1'b0,io_b[479 : 432]});
  assign _zz__zz_io_s_27_2 = _zz_io_s_26;
  assign _zz__zz_io_s_27_1 = {48'd0, _zz__zz_io_s_27_2};
  assign _zz__zz_io_s_30 = ({1'b0,io_a[527 : 480]} + {1'b0,io_b[527 : 480]});
  assign _zz__zz_io_s_30_2 = _zz_io_s_29;
  assign _zz__zz_io_s_30_1 = {48'd0, _zz__zz_io_s_30_2};
  assign _zz__zz_io_s_33 = ({1'b0,io_a[575 : 528]} + {1'b0,io_b[575 : 528]});
  assign _zz__zz_io_s_33_2 = _zz_io_s_32;
  assign _zz__zz_io_s_33_1 = {48'd0, _zz__zz_io_s_33_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[239 : 192] = _zz_io_s_13;
    io_s[287 : 240] = _zz_io_s_16;
    io_s[335 : 288] = _zz_io_s_19;
    io_s[383 : 336] = _zz_io_s_22;
    io_s[431 : 384] = _zz_io_s_25;
    io_s[479 : 432] = _zz_io_s_28;
    io_s[527 : 480] = _zz_io_s_31;
    io_s[575 : 528] = _zz_io_s_34;
    io_s[576] = _zz_io_s_36;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_1);
  assign _zz_io_s_18 = (_zz__zz_io_s_18 + _zz__zz_io_s_18_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  assign _zz_io_s_24 = (_zz__zz_io_s_24 + _zz__zz_io_s_24_1);
  assign _zz_io_s_27 = (_zz__zz_io_s_27 + _zz__zz_io_s_27_1);
  assign _zz_io_s_30 = (_zz__zz_io_s_30 + _zz__zz_io_s_30_1);
  assign _zz_io_s_33 = (_zz__zz_io_s_33 + _zz__zz_io_s_33_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_13 <= _zz_io_s_12[47:0];
    _zz_io_s_14 <= _zz_io_s_12[48];
    _zz_io_s_16 <= _zz_io_s_15[47:0];
    _zz_io_s_17 <= _zz_io_s_15[48];
    _zz_io_s_19 <= _zz_io_s_18[47:0];
    _zz_io_s_20 <= _zz_io_s_18[48];
    _zz_io_s_22 <= _zz_io_s_21[47:0];
    _zz_io_s_23 <= _zz_io_s_21[48];
    _zz_io_s_25 <= _zz_io_s_24[47:0];
    _zz_io_s_26 <= _zz_io_s_24[48];
    _zz_io_s_28 <= _zz_io_s_27[47:0];
    _zz_io_s_29 <= _zz_io_s_27[48];
    _zz_io_s_31 <= _zz_io_s_30[47:0];
    _zz_io_s_32 <= _zz_io_s_30[48];
    _zz_io_s_34 <= _zz_io_s_33[47:0];
    _zz_io_s_35 <= _zz_io_s_33[48];
    _zz_io_s_36 <= _zz_io_s_35;
  end


endmodule

module BADD_655 (
  input      [384:0]  io_a,
  input      [384:0]  io_b,
  input               io_c,
  output reg [385:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [384:0]  _zz__zz_io_s_1;
  wire       [48:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [384:0]  _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_3_3;
  wire       [0:0]    _zz__zz_io_s_3_4;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [384:0]  _zz__zz_io_s_6_1;
  wire       [48:0]   _zz__zz_io_s_6_2;
  wire       [0:0]    _zz__zz_io_s_6_3;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [384:0]  _zz__zz_io_s_9_1;
  wire       [48:0]   _zz__zz_io_s_9_2;
  wire       [0:0]    _zz__zz_io_s_9_3;
  wire       [48:0]   _zz__zz_io_s_12;
  wire       [384:0]  _zz__zz_io_s_12_1;
  wire       [48:0]   _zz__zz_io_s_12_2;
  wire       [0:0]    _zz__zz_io_s_12_3;
  wire       [48:0]   _zz__zz_io_s_15;
  wire       [384:0]  _zz__zz_io_s_15_1;
  wire       [48:0]   _zz__zz_io_s_15_2;
  wire       [0:0]    _zz__zz_io_s_15_3;
  wire       [48:0]   _zz__zz_io_s_18;
  wire       [384:0]  _zz__zz_io_s_18_1;
  wire       [48:0]   _zz__zz_io_s_18_2;
  wire       [0:0]    _zz__zz_io_s_18_3;
  wire       [48:0]   _zz__zz_io_s_21;
  wire       [384:0]  _zz__zz_io_s_21_1;
  wire       [48:0]   _zz__zz_io_s_21_2;
  wire       [0:0]    _zz__zz_io_s_21_3;
  wire       [1:0]    _zz__zz_io_s_24;
  wire       [384:0]  _zz__zz_io_s_24_1;
  wire       [1:0]    _zz__zz_io_s_24_2;
  wire       [0:0]    _zz__zz_io_s_24_3;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [48:0]   _zz_io_s_12;
  reg        [47:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [48:0]   _zz_io_s_15;
  reg        [47:0]   _zz_io_s_16;
  reg                 _zz_io_s_17;
  wire       [48:0]   _zz_io_s_18;
  reg        [47:0]   _zz_io_s_19;
  reg                 _zz_io_s_20;
  wire       [48:0]   _zz_io_s_21;
  reg        [47:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  wire       [1:0]    _zz_io_s_24;
  reg        [0:0]    _zz_io_s_25;
  reg                 _zz_io_s_26;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,_zz__zz_io_s_1[47 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {48'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_3_1 = ({1'b0,io_a[95 : 48]} + {1'b0,_zz__zz_io_s_3_2[95 : 48]});
  assign _zz__zz_io_s_3_2 = (~ io_b);
  assign _zz__zz_io_s_3_4 = _zz_io_s_2;
  assign _zz__zz_io_s_3_3 = {48'd0, _zz__zz_io_s_3_4};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,_zz__zz_io_s_6_1[143 : 96]});
  assign _zz__zz_io_s_6_1 = (~ io_b);
  assign _zz__zz_io_s_6_3 = _zz_io_s_5;
  assign _zz__zz_io_s_6_2 = {48'd0, _zz__zz_io_s_6_3};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,_zz__zz_io_s_9_1[191 : 144]});
  assign _zz__zz_io_s_9_1 = (~ io_b);
  assign _zz__zz_io_s_9_3 = _zz_io_s_8;
  assign _zz__zz_io_s_9_2 = {48'd0, _zz__zz_io_s_9_3};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[239 : 192]} + {1'b0,_zz__zz_io_s_12_1[239 : 192]});
  assign _zz__zz_io_s_12_1 = (~ io_b);
  assign _zz__zz_io_s_12_3 = _zz_io_s_11;
  assign _zz__zz_io_s_12_2 = {48'd0, _zz__zz_io_s_12_3};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[287 : 240]} + {1'b0,_zz__zz_io_s_15_1[287 : 240]});
  assign _zz__zz_io_s_15_1 = (~ io_b);
  assign _zz__zz_io_s_15_3 = _zz_io_s_14;
  assign _zz__zz_io_s_15_2 = {48'd0, _zz__zz_io_s_15_3};
  assign _zz__zz_io_s_18 = ({1'b0,io_a[335 : 288]} + {1'b0,_zz__zz_io_s_18_1[335 : 288]});
  assign _zz__zz_io_s_18_1 = (~ io_b);
  assign _zz__zz_io_s_18_3 = _zz_io_s_17;
  assign _zz__zz_io_s_18_2 = {48'd0, _zz__zz_io_s_18_3};
  assign _zz__zz_io_s_21 = ({1'b0,io_a[383 : 336]} + {1'b0,_zz__zz_io_s_21_1[383 : 336]});
  assign _zz__zz_io_s_21_1 = (~ io_b);
  assign _zz__zz_io_s_21_3 = _zz_io_s_20;
  assign _zz__zz_io_s_21_2 = {48'd0, _zz__zz_io_s_21_3};
  assign _zz__zz_io_s_24 = ({1'b0,io_a[384 : 384]} + {1'b0,_zz__zz_io_s_24_1[384 : 384]});
  assign _zz__zz_io_s_24_1 = (~ io_b);
  assign _zz__zz_io_s_24_3 = _zz_io_s_23;
  assign _zz__zz_io_s_24_2 = {1'd0, _zz__zz_io_s_24_3};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[239 : 192] = _zz_io_s_13;
    io_s[287 : 240] = _zz_io_s_16;
    io_s[335 : 288] = _zz_io_s_19;
    io_s[383 : 336] = _zz_io_s_22;
    io_s[384 : 384] = _zz_io_s_25;
    io_s[385] = (! _zz_io_s_26);
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3_1 + _zz__zz_io_s_3_3);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_2);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_2);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_2);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_2);
  assign _zz_io_s_18 = (_zz__zz_io_s_18 + _zz__zz_io_s_18_2);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_2);
  assign _zz_io_s_24 = (_zz__zz_io_s_24 + _zz__zz_io_s_24_2);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_13 <= _zz_io_s_12[47:0];
    _zz_io_s_14 <= _zz_io_s_12[48];
    _zz_io_s_16 <= _zz_io_s_15[47:0];
    _zz_io_s_17 <= _zz_io_s_15[48];
    _zz_io_s_19 <= _zz_io_s_18[47:0];
    _zz_io_s_20 <= _zz_io_s_18[48];
    _zz_io_s_22 <= _zz_io_s_21[47:0];
    _zz_io_s_23 <= _zz_io_s_21[48];
    _zz_io_s_25 <= _zz_io_s_24[0:0];
    _zz_io_s_26 <= _zz_io_s_24[1];
  end


endmodule

module BADD_654 (
  input      [383:0]  io_a,
  input      [383:0]  io_b,
  input               io_c,
  output reg [384:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [48:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [48:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [48:0]   _zz__zz_io_s_12;
  wire       [48:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [48:0]   _zz__zz_io_s_15;
  wire       [48:0]   _zz__zz_io_s_15_1;
  wire       [0:0]    _zz__zz_io_s_15_2;
  wire       [48:0]   _zz__zz_io_s_18;
  wire       [48:0]   _zz__zz_io_s_18_1;
  wire       [0:0]    _zz__zz_io_s_18_2;
  wire       [48:0]   _zz__zz_io_s_21;
  wire       [48:0]   _zz__zz_io_s_21_1;
  wire       [0:0]    _zz__zz_io_s_21_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [48:0]   _zz_io_s_12;
  reg        [47:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [48:0]   _zz_io_s_15;
  reg        [47:0]   _zz_io_s_16;
  reg                 _zz_io_s_17;
  wire       [48:0]   _zz_io_s_18;
  reg        [47:0]   _zz_io_s_19;
  reg                 _zz_io_s_20;
  wire       [48:0]   _zz_io_s_21;
  reg        [47:0]   _zz_io_s_22;
  reg                 _zz_io_s_23;
  reg                 _zz_io_s_24;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,io_b[143 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {48'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,io_b[191 : 144]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {48'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[239 : 192]} + {1'b0,io_b[239 : 192]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {48'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[287 : 240]} + {1'b0,io_b[287 : 240]});
  assign _zz__zz_io_s_15_2 = _zz_io_s_14;
  assign _zz__zz_io_s_15_1 = {48'd0, _zz__zz_io_s_15_2};
  assign _zz__zz_io_s_18 = ({1'b0,io_a[335 : 288]} + {1'b0,io_b[335 : 288]});
  assign _zz__zz_io_s_18_2 = _zz_io_s_17;
  assign _zz__zz_io_s_18_1 = {48'd0, _zz__zz_io_s_18_2};
  assign _zz__zz_io_s_21 = ({1'b0,io_a[383 : 336]} + {1'b0,io_b[383 : 336]});
  assign _zz__zz_io_s_21_2 = _zz_io_s_20;
  assign _zz__zz_io_s_21_1 = {48'd0, _zz__zz_io_s_21_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[239 : 192] = _zz_io_s_13;
    io_s[287 : 240] = _zz_io_s_16;
    io_s[335 : 288] = _zz_io_s_19;
    io_s[383 : 336] = _zz_io_s_22;
    io_s[384] = _zz_io_s_24;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_1);
  assign _zz_io_s_18 = (_zz__zz_io_s_18 + _zz__zz_io_s_18_1);
  assign _zz_io_s_21 = (_zz__zz_io_s_21 + _zz__zz_io_s_21_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_13 <= _zz_io_s_12[47:0];
    _zz_io_s_14 <= _zz_io_s_12[48];
    _zz_io_s_16 <= _zz_io_s_15[47:0];
    _zz_io_s_17 <= _zz_io_s_15[48];
    _zz_io_s_19 <= _zz_io_s_18[47:0];
    _zz_io_s_20 <= _zz_io_s_18[48];
    _zz_io_s_22 <= _zz_io_s_21[47:0];
    _zz_io_s_23 <= _zz_io_s_21[48];
    _zz_io_s_24 <= _zz_io_s_23;
  end


endmodule

module KaratsubaCore_71 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_a_2,
  input      [47:0]   io_a_3,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  input      [47:0]   io_b_2,
  input      [47:0]   io_b_3,
  output reg [383:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [192:0]  karatsuba_add2_io_a;
  wire       [287:0]  karatsuba_noExtend_add3_io_a;
  reg        [287:0]  karatsuba_noExtend_add3_io_b;
  wire       [191:0]  karatsuba_lsbMul_io_p;
  wire       [193:0]  karatsuba_midMul_io_p;
  wire       [191:0]  karatsuba_msbMul_io_p;
  wire       [192:0]  karatsuba_add1_io_s;
  wire       [193:0]  karatsuba_add2_io_s;
  wire       [288:0]  karatsuba_noExtend_add3_io_s;
  wire       [192:0]  _zz_io_a;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_a_1;
  reg        [48:0]   _zz_io_b_0;
  reg        [48:0]   _zz_io_b_1;
  reg        [192:0]  karatsuba_msbMul_karatsuba_add1_io_s_delay_1;
  reg        [95:0]   _zz_io_b;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4;
  reg        [191:0]  karatsuba_msbMul_karatsuba_msbMul_io_p_delay_5;
  reg        [95:0]   _zz_io_p;
  reg        [95:0]   _zz_io_p_1;

  assign _zz_io_a = karatsuba_add2_io_s[192:0];
  KaratsubaCore_231 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]                ), //i
    .io_a_1 (io_a_1[47:0]                ), //i
    .io_b_0 (io_b_0[47:0]                ), //i
    .io_b_1 (io_b_1[47:0]                ), //i
    .io_p   (karatsuba_lsbMul_io_p[191:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_232 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]            ), //i
    .io_a_1 (_zz_io_a_1[48:0]            ), //i
    .io_b_0 (_zz_io_b_0[48:0]            ), //i
    .io_b_1 (_zz_io_b_1[48:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[193:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_233 karatsuba_msbMul (
    .io_a_0 (io_a_2[47:0]                ), //i
    .io_a_1 (io_a_3[47:0]                ), //i
    .io_b_0 (io_b_2[47:0]                ), //i
    .io_b_1 (io_b_3[47:0]                ), //i
    .io_p   (karatsuba_msbMul_io_p[191:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_834 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[191:0]), //i
    .io_b   (karatsuba_msbMul_io_p[191:0]), //i
    .io_c   (1'b0                        ), //i
    .io_s   (karatsuba_add1_io_s[192:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_835 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[192:0]                         ), //i
    .io_b   (karatsuba_msbMul_karatsuba_add1_io_s_delay_1[192:0]), //i
    .io_c   (1'b1                                               ), //i
    .io_s   (karatsuba_add2_io_s[193:0]                         ), //o
    .clk    (clk                                                ), //i
    .resetn (resetn                                             )  //i
  );
  BADD_836 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[287:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[287:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[288:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[192:0];
  assign karatsuba_noExtend_add3_io_a = {95'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[95 : 0] = _zz_io_b;
    karatsuba_noExtend_add3_io_b[287 : 96] = karatsuba_msbMul_karatsuba_msbMul_io_p_delay_5;
  end

  always @(*) begin
    io_p[95 : 0] = _zz_io_p_1;
    io_p[383 : 96] = karatsuba_noExtend_add3_io_s[287:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_2});
    _zz_io_a_1 <= ({1'b0,io_a_1} + {1'b0,io_a_3});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_2});
    _zz_io_b_1 <= ({1'b0,io_b_1} + {1'b0,io_b_3});
    karatsuba_msbMul_karatsuba_add1_io_s_delay_1 <= karatsuba_add1_io_s;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 96);
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_5 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4;
    _zz_io_p <= karatsuba_lsbMul_io_p[95 : 0];
    _zz_io_p_1 <= _zz_io_p;
  end


endmodule

module KaratsubaCore_70 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_a_1,
  input      [48:0]   io_a_2,
  input      [48:0]   io_a_3,
  input      [48:0]   io_b_0,
  input      [48:0]   io_b_1,
  input      [48:0]   io_b_2,
  input      [48:0]   io_b_3,
  output reg [385:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [194:0]  karatsuba_add2_io_a;
  wire       [194:0]  karatsuba_hasExtend_add3_io_a;
  wire       [194:0]  karatsuba_hasExtend_add3_io_b;
  wire       [193:0]  karatsuba_hasExtend_add4_io_a;
  wire       [193:0]  karatsuba_lsbMul_io_p;
  wire       [195:0]  karatsuba_midMul_io_p;
  wire       [193:0]  karatsuba_msbMul_io_p;
  wire       [194:0]  karatsuba_add1_io_s;
  wire       [195:0]  karatsuba_add2_io_s;
  wire       [195:0]  karatsuba_hasExtend_add3_io_s;
  wire       [194:0]  karatsuba_hasExtend_add4_io_s;
  wire       [97:0]   _zz_io_b;
  wire       [99:0]   _zz_io_a;
  reg        [49:0]   _zz_io_a_0;
  reg        [49:0]   _zz_io_a_1;
  reg        [49:0]   _zz_io_b_0;
  reg        [49:0]   _zz_io_b_1;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_4;
  reg        [193:0]  karatsuba_midMul_karatsuba_msbMul_io_p_delay_5;
  reg        [95:0]   _zz_io_p;
  reg        [95:0]   _zz_io_p_1;
  reg        [95:0]   _zz_io_p_2;

  assign _zz_io_b = (karatsuba_lsbMul_io_p >>> 96);
  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 96);
  KaratsubaCore_228 karatsuba_lsbMul (
    .io_a_0 (io_a_0[48:0]                ), //i
    .io_a_1 (io_a_1[48:0]                ), //i
    .io_b_0 (io_b_0[48:0]                ), //i
    .io_b_1 (io_b_1[48:0]                ), //i
    .io_p   (karatsuba_lsbMul_io_p[193:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_229 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[49:0]            ), //i
    .io_a_1 (_zz_io_a_1[49:0]            ), //i
    .io_b_0 (_zz_io_b_0[49:0]            ), //i
    .io_b_1 (_zz_io_b_1[49:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[195:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_230 karatsuba_msbMul (
    .io_a_0 (io_a_2[48:0]                ), //i
    .io_a_1 (io_a_3[48:0]                ), //i
    .io_b_0 (io_b_2[48:0]                ), //i
    .io_b_1 (io_b_3[48:0]                ), //i
    .io_p   (karatsuba_msbMul_io_p[193:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_830 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[193:0]), //i
    .io_b   (karatsuba_msbMul_io_p[193:0]), //i
    .io_c   (1'b0                        ), //i
    .io_s   (karatsuba_add1_io_s[194:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_831 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[194:0]), //i
    .io_b   (karatsuba_add1_io_s[194:0]), //i
    .io_c   (1'b1                      ), //i
    .io_s   (karatsuba_add2_io_s[195:0]), //o
    .clk    (clk                       ), //i
    .resetn (resetn                    )  //i
  );
  BADD_832 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[194:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[194:0]), //i
    .io_c   (1'b0                                ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[195:0]), //o
    .clk    (clk                                 ), //i
    .resetn (resetn                              )  //i
  );
  BADD_830 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[193:0]                 ), //i
    .io_b   (karatsuba_midMul_karatsuba_msbMul_io_p_delay_5[193:0]), //i
    .io_c   (1'b0                                                 ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[194:0]                 ), //o
    .clk    (clk                                                  ), //i
    .resetn (resetn                                               )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[194:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[194:0];
  assign karatsuba_hasExtend_add3_io_b = {97'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {94'd0, _zz_io_a};
  always @(*) begin
    io_p[95 : 0] = _zz_io_p_1;
    io_p[191 : 96] = _zz_io_p_2;
    io_p[385 : 192] = karatsuba_hasExtend_add4_io_s[193:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_2});
    _zz_io_a_1 <= ({1'b0,io_a_1} + {1'b0,io_a_3});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_2});
    _zz_io_b_1 <= ({1'b0,io_b_1} + {1'b0,io_b_3});
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_5 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_4;
    _zz_io_p <= karatsuba_lsbMul_io_p[95 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= karatsuba_hasExtend_add3_io_s[95:0];
  end


endmodule

module KaratsubaCore_69 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_a_2,
  input      [47:0]   io_a_3,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  input      [47:0]   io_b_2,
  input      [47:0]   io_b_3,
  output reg [383:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [192:0]  karatsuba_add2_io_a;
  wire       [287:0]  karatsuba_noExtend_add3_io_a;
  reg        [287:0]  karatsuba_noExtend_add3_io_b;
  wire       [191:0]  karatsuba_lsbMul_io_p;
  wire       [193:0]  karatsuba_midMul_io_p;
  wire       [191:0]  karatsuba_msbMul_io_p;
  wire       [192:0]  karatsuba_add1_io_s;
  wire       [193:0]  karatsuba_add2_io_s;
  wire       [288:0]  karatsuba_noExtend_add3_io_s;
  wire       [192:0]  _zz_io_a;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_a_1;
  reg        [48:0]   _zz_io_b_0;
  reg        [48:0]   _zz_io_b_1;
  reg        [192:0]  karatsuba_lsbMul_karatsuba_add1_io_s_delay_1;
  reg        [95:0]   _zz_io_b;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4;
  reg        [191:0]  karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_5;
  reg        [95:0]   _zz_io_p;
  reg        [95:0]   _zz_io_p_1;

  assign _zz_io_a = karatsuba_add2_io_s[192:0];
  KaratsubaCore_231 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]                ), //i
    .io_a_1 (io_a_1[47:0]                ), //i
    .io_b_0 (io_b_0[47:0]                ), //i
    .io_b_1 (io_b_1[47:0]                ), //i
    .io_p   (karatsuba_lsbMul_io_p[191:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_232 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]            ), //i
    .io_a_1 (_zz_io_a_1[48:0]            ), //i
    .io_b_0 (_zz_io_b_0[48:0]            ), //i
    .io_b_1 (_zz_io_b_1[48:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[193:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_233 karatsuba_msbMul (
    .io_a_0 (io_a_2[47:0]                ), //i
    .io_a_1 (io_a_3[47:0]                ), //i
    .io_b_0 (io_b_2[47:0]                ), //i
    .io_b_1 (io_b_3[47:0]                ), //i
    .io_p   (karatsuba_msbMul_io_p[191:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_834 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[191:0]), //i
    .io_b   (karatsuba_msbMul_io_p[191:0]), //i
    .io_c   (1'b0                        ), //i
    .io_s   (karatsuba_add1_io_s[192:0]  ), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  BADD_835 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[192:0]                         ), //i
    .io_b   (karatsuba_lsbMul_karatsuba_add1_io_s_delay_1[192:0]), //i
    .io_c   (1'b1                                               ), //i
    .io_s   (karatsuba_add2_io_s[193:0]                         ), //o
    .clk    (clk                                                ), //i
    .resetn (resetn                                             )  //i
  );
  BADD_836 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[287:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[287:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[288:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[192:0];
  assign karatsuba_noExtend_add3_io_a = {95'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[95 : 0] = _zz_io_b;
    karatsuba_noExtend_add3_io_b[287 : 96] = karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_5;
  end

  always @(*) begin
    io_p[95 : 0] = _zz_io_p_1;
    io_p[383 : 96] = karatsuba_noExtend_add3_io_s[287:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_2});
    _zz_io_a_1 <= ({1'b0,io_a_1} + {1'b0,io_a_3});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_2});
    _zz_io_b_1 <= ({1'b0,io_b_1} + {1'b0,io_b_3});
    karatsuba_lsbMul_karatsuba_add1_io_s_delay_1 <= karatsuba_add1_io_s;
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 96);
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_5 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4;
    _zz_io_p <= karatsuba_lsbMul_io_p[95 : 0];
    _zz_io_p_1 <= _zz_io_p;
  end


endmodule

//BADD_659 replaced by BADD_836

//BADD_658 replaced by BADD_835

//BADD_657 replaced by BADD_834

//KaratsubaCore_74 replaced by KaratsubaCore_233

//KaratsubaCore_73 replaced by KaratsubaCore_232

//KaratsubaCore_72 replaced by KaratsubaCore_231

//BADD_663 replaced by BADD_830

//BADD_662 replaced by BADD_832

//BADD_661 replaced by BADD_831

//BADD_660 replaced by BADD_830

//KaratsubaCore_77 replaced by KaratsubaCore_230

//KaratsubaCore_76 replaced by KaratsubaCore_229

//KaratsubaCore_75 replaced by KaratsubaCore_228

//BADD_666 replaced by BADD_836

//BADD_665 replaced by BADD_835

//BADD_664 replaced by BADD_834

//KaratsubaCore_80 replaced by KaratsubaCore_233

//KaratsubaCore_79 replaced by KaratsubaCore_232

//KaratsubaCore_78 replaced by KaratsubaCore_231

//BADD_669 replaced by BADD_836

//BADD_668 replaced by BADD_835

//BADD_667 replaced by BADD_834

//KaratsubaCore_83 replaced by KaratsubaCore_233

//KaratsubaCore_82 replaced by KaratsubaCore_232

//KaratsubaCore_81 replaced by KaratsubaCore_231

//BADD_673 replaced by BADD_830

//BADD_672 replaced by BADD_832

//BADD_671 replaced by BADD_831

//BADD_670 replaced by BADD_830

//KaratsubaCore_86 replaced by KaratsubaCore_230

//KaratsubaCore_85 replaced by KaratsubaCore_229

//KaratsubaCore_84 replaced by KaratsubaCore_228

//BADD_676 replaced by BADD_836

//BADD_675 replaced by BADD_835

//BADD_674 replaced by BADD_834

//KaratsubaCore_89 replaced by KaratsubaCore_233

//KaratsubaCore_88 replaced by KaratsubaCore_232

//KaratsubaCore_87 replaced by KaratsubaCore_231

//BADD_679 replaced by BADD_836

//BADD_678 replaced by BADD_835

//BADD_677 replaced by BADD_834

//KaratsubaCore_92 replaced by KaratsubaCore_233

//KaratsubaCore_91 replaced by KaratsubaCore_232

//KaratsubaCore_90 replaced by KaratsubaCore_231

//BADD_683 replaced by BADD_830

//BADD_682 replaced by BADD_832

//BADD_681 replaced by BADD_831

//BADD_680 replaced by BADD_830

//KaratsubaCore_95 replaced by KaratsubaCore_230

//KaratsubaCore_94 replaced by KaratsubaCore_229

//KaratsubaCore_93 replaced by KaratsubaCore_228

//BADD_686 replaced by BADD_836

//BADD_685 replaced by BADD_835

//BADD_684 replaced by BADD_834

//KaratsubaCore_98 replaced by KaratsubaCore_233

//KaratsubaCore_97 replaced by KaratsubaCore_232

//KaratsubaCore_96 replaced by KaratsubaCore_231

//BADD_689 replaced by BADD_836

//BADD_688 replaced by BADD_835

//BADD_687 replaced by BADD_834

//KaratsubaCore_101 replaced by KaratsubaCore_233

//KaratsubaCore_100 replaced by KaratsubaCore_232

//KaratsubaCore_99 replaced by KaratsubaCore_231

//BADD_693 replaced by BADD_830

//BADD_692 replaced by BADD_832

//BADD_691 replaced by BADD_831

//BADD_690 replaced by BADD_830

//KaratsubaCore_104 replaced by KaratsubaCore_230

//KaratsubaCore_103 replaced by KaratsubaCore_229

//KaratsubaCore_102 replaced by KaratsubaCore_228

//BADD_696 replaced by BADD_836

//BADD_695 replaced by BADD_835

//BADD_694 replaced by BADD_834

//KaratsubaCore_107 replaced by KaratsubaCore_233

//KaratsubaCore_106 replaced by KaratsubaCore_232

//KaratsubaCore_105 replaced by KaratsubaCore_231

//BADD_699 replaced by BADD_836

//BADD_698 replaced by BADD_835

//BADD_697 replaced by BADD_834

//KaratsubaCore_110 replaced by KaratsubaCore_233

//KaratsubaCore_109 replaced by KaratsubaCore_232

//KaratsubaCore_108 replaced by KaratsubaCore_231

//BADD_703 replaced by BADD_830

//BADD_702 replaced by BADD_832

//BADD_701 replaced by BADD_831

//BADD_700 replaced by BADD_830

//KaratsubaCore_113 replaced by KaratsubaCore_230

//KaratsubaCore_112 replaced by KaratsubaCore_229

//KaratsubaCore_111 replaced by KaratsubaCore_228

//BADD_706 replaced by BADD_836

//BADD_705 replaced by BADD_835

//BADD_704 replaced by BADD_834

//KaratsubaCore_116 replaced by KaratsubaCore_233

//KaratsubaCore_115 replaced by KaratsubaCore_232

//KaratsubaCore_114 replaced by KaratsubaCore_231

//BADD_709 replaced by BADD_836

//BADD_708 replaced by BADD_835

//BADD_707 replaced by BADD_834

//KaratsubaCore_119 replaced by KaratsubaCore_233

//KaratsubaCore_118 replaced by KaratsubaCore_232

//KaratsubaCore_117 replaced by KaratsubaCore_231

//BADD_713 replaced by BADD_830

//BADD_712 replaced by BADD_832

//BADD_711 replaced by BADD_831

//BADD_710 replaced by BADD_830

//KaratsubaCore_122 replaced by KaratsubaCore_230

//KaratsubaCore_121 replaced by KaratsubaCore_229

//KaratsubaCore_120 replaced by KaratsubaCore_228

//BADD_716 replaced by BADD_836

//BADD_715 replaced by BADD_835

//BADD_714 replaced by BADD_834

//KaratsubaCore_125 replaced by KaratsubaCore_233

//KaratsubaCore_124 replaced by KaratsubaCore_232

//KaratsubaCore_123 replaced by KaratsubaCore_231

//BADD_719 replaced by BADD_836

//BADD_718 replaced by BADD_835

//BADD_717 replaced by BADD_834

//KaratsubaCore_128 replaced by KaratsubaCore_233

//KaratsubaCore_127 replaced by KaratsubaCore_232

//KaratsubaCore_126 replaced by KaratsubaCore_231

//BADD_723 replaced by BADD_830

//BADD_722 replaced by BADD_832

//BADD_721 replaced by BADD_831

//BADD_720 replaced by BADD_830

//KaratsubaCore_131 replaced by KaratsubaCore_230

//KaratsubaCore_130 replaced by KaratsubaCore_229

//KaratsubaCore_129 replaced by KaratsubaCore_228

//BADD_726 replaced by BADD_836

//BADD_725 replaced by BADD_835

//BADD_724 replaced by BADD_834

//KaratsubaCore_134 replaced by KaratsubaCore_233

//KaratsubaCore_133 replaced by KaratsubaCore_232

//KaratsubaCore_132 replaced by KaratsubaCore_231

//BADD_729 replaced by BADD_836

//BADD_728 replaced by BADD_835

//BADD_727 replaced by BADD_834

//KaratsubaCore_137 replaced by KaratsubaCore_233

//KaratsubaCore_136 replaced by KaratsubaCore_232

//KaratsubaCore_135 replaced by KaratsubaCore_231

//BADD_733 replaced by BADD_830

//BADD_732 replaced by BADD_832

//BADD_731 replaced by BADD_831

//BADD_730 replaced by BADD_830

//KaratsubaCore_140 replaced by KaratsubaCore_230

//KaratsubaCore_139 replaced by KaratsubaCore_229

//KaratsubaCore_138 replaced by KaratsubaCore_228

//BADD_736 replaced by BADD_836

//BADD_735 replaced by BADD_835

//BADD_734 replaced by BADD_834

//KaratsubaCore_143 replaced by KaratsubaCore_233

//KaratsubaCore_142 replaced by KaratsubaCore_232

//KaratsubaCore_141 replaced by KaratsubaCore_231

//BADD_739 replaced by BADD_836

//BADD_738 replaced by BADD_835

//BADD_737 replaced by BADD_834

//KaratsubaCore_146 replaced by KaratsubaCore_233

//KaratsubaCore_145 replaced by KaratsubaCore_232

//KaratsubaCore_144 replaced by KaratsubaCore_231

//BADD_743 replaced by BADD_830

//BADD_742 replaced by BADD_832

//BADD_741 replaced by BADD_831

//BADD_740 replaced by BADD_830

//KaratsubaCore_149 replaced by KaratsubaCore_230

//KaratsubaCore_148 replaced by KaratsubaCore_229

//KaratsubaCore_147 replaced by KaratsubaCore_228

//BADD_746 replaced by BADD_836

//BADD_745 replaced by BADD_835

//BADD_744 replaced by BADD_834

//KaratsubaCore_152 replaced by KaratsubaCore_233

//KaratsubaCore_151 replaced by KaratsubaCore_232

//KaratsubaCore_150 replaced by KaratsubaCore_231

//BADD_749 replaced by BADD_836

//BADD_748 replaced by BADD_835

//BADD_747 replaced by BADD_834

//KaratsubaCore_155 replaced by KaratsubaCore_233

//KaratsubaCore_154 replaced by KaratsubaCore_232

//KaratsubaCore_153 replaced by KaratsubaCore_231

//BADD_753 replaced by BADD_830

//BADD_752 replaced by BADD_832

//BADD_751 replaced by BADD_831

//BADD_750 replaced by BADD_830

//KaratsubaCore_158 replaced by KaratsubaCore_230

//KaratsubaCore_157 replaced by KaratsubaCore_229

//KaratsubaCore_156 replaced by KaratsubaCore_228

//BADD_756 replaced by BADD_836

//BADD_755 replaced by BADD_835

//BADD_754 replaced by BADD_834

//KaratsubaCore_161 replaced by KaratsubaCore_233

//KaratsubaCore_160 replaced by KaratsubaCore_232

//KaratsubaCore_159 replaced by KaratsubaCore_231

//BADD_759 replaced by BADD_836

//BADD_758 replaced by BADD_835

//BADD_757 replaced by BADD_834

//KaratsubaCore_164 replaced by KaratsubaCore_233

//KaratsubaCore_163 replaced by KaratsubaCore_232

//KaratsubaCore_162 replaced by KaratsubaCore_231

//BADD_763 replaced by BADD_830

//BADD_762 replaced by BADD_832

//BADD_761 replaced by BADD_831

//BADD_760 replaced by BADD_830

//KaratsubaCore_167 replaced by KaratsubaCore_230

//KaratsubaCore_166 replaced by KaratsubaCore_229

//KaratsubaCore_165 replaced by KaratsubaCore_228

//BADD_766 replaced by BADD_836

//BADD_765 replaced by BADD_835

//BADD_764 replaced by BADD_834

//KaratsubaCore_170 replaced by KaratsubaCore_233

//KaratsubaCore_169 replaced by KaratsubaCore_232

//KaratsubaCore_168 replaced by KaratsubaCore_231

//BADD_769 replaced by BADD_836

//BADD_768 replaced by BADD_835

//BADD_767 replaced by BADD_834

//KaratsubaCore_173 replaced by KaratsubaCore_233

//KaratsubaCore_172 replaced by KaratsubaCore_232

//KaratsubaCore_171 replaced by KaratsubaCore_231

//BADD_773 replaced by BADD_830

//BADD_772 replaced by BADD_832

//BADD_771 replaced by BADD_831

//BADD_770 replaced by BADD_830

//KaratsubaCore_176 replaced by KaratsubaCore_230

//KaratsubaCore_175 replaced by KaratsubaCore_229

//KaratsubaCore_174 replaced by KaratsubaCore_228

//BADD_776 replaced by BADD_836

//BADD_775 replaced by BADD_835

//BADD_774 replaced by BADD_834

//KaratsubaCore_179 replaced by KaratsubaCore_233

//KaratsubaCore_178 replaced by KaratsubaCore_232

//KaratsubaCore_177 replaced by KaratsubaCore_231

//BADD_779 replaced by BADD_836

//BADD_778 replaced by BADD_835

//BADD_777 replaced by BADD_834

//KaratsubaCore_182 replaced by KaratsubaCore_233

//KaratsubaCore_181 replaced by KaratsubaCore_232

//KaratsubaCore_180 replaced by KaratsubaCore_231

//BADD_783 replaced by BADD_830

//BADD_782 replaced by BADD_832

//BADD_781 replaced by BADD_831

//BADD_780 replaced by BADD_830

//KaratsubaCore_185 replaced by KaratsubaCore_230

//KaratsubaCore_184 replaced by KaratsubaCore_229

//KaratsubaCore_183 replaced by KaratsubaCore_228

//BADD_786 replaced by BADD_836

//BADD_785 replaced by BADD_835

//BADD_784 replaced by BADD_834

//KaratsubaCore_188 replaced by KaratsubaCore_233

//KaratsubaCore_187 replaced by KaratsubaCore_232

//KaratsubaCore_186 replaced by KaratsubaCore_231

//BADD_789 replaced by BADD_836

//BADD_788 replaced by BADD_835

//BADD_787 replaced by BADD_834

//KaratsubaCore_191 replaced by KaratsubaCore_233

//KaratsubaCore_190 replaced by KaratsubaCore_232

//KaratsubaCore_189 replaced by KaratsubaCore_231

//BADD_793 replaced by BADD_830

//BADD_792 replaced by BADD_832

//BADD_791 replaced by BADD_831

//BADD_790 replaced by BADD_830

//KaratsubaCore_194 replaced by KaratsubaCore_230

//KaratsubaCore_193 replaced by KaratsubaCore_229

//KaratsubaCore_192 replaced by KaratsubaCore_228

//BADD_796 replaced by BADD_836

//BADD_795 replaced by BADD_835

//BADD_794 replaced by BADD_834

//KaratsubaCore_197 replaced by KaratsubaCore_233

//KaratsubaCore_196 replaced by KaratsubaCore_232

//KaratsubaCore_195 replaced by KaratsubaCore_231

//BADD_799 replaced by BADD_836

//BADD_798 replaced by BADD_835

//BADD_797 replaced by BADD_834

//KaratsubaCore_200 replaced by KaratsubaCore_233

//KaratsubaCore_199 replaced by KaratsubaCore_232

//KaratsubaCore_198 replaced by KaratsubaCore_231

//BADD_803 replaced by BADD_830

//BADD_802 replaced by BADD_832

//BADD_801 replaced by BADD_831

//BADD_800 replaced by BADD_830

//KaratsubaCore_203 replaced by KaratsubaCore_230

//KaratsubaCore_202 replaced by KaratsubaCore_229

//KaratsubaCore_201 replaced by KaratsubaCore_228

//BADD_806 replaced by BADD_836

//BADD_805 replaced by BADD_835

//BADD_804 replaced by BADD_834

//KaratsubaCore_206 replaced by KaratsubaCore_233

//KaratsubaCore_205 replaced by KaratsubaCore_232

//KaratsubaCore_204 replaced by KaratsubaCore_231

//BADD_809 replaced by BADD_836

//BADD_808 replaced by BADD_835

//BADD_807 replaced by BADD_834

//KaratsubaCore_209 replaced by KaratsubaCore_233

//KaratsubaCore_208 replaced by KaratsubaCore_232

//KaratsubaCore_207 replaced by KaratsubaCore_231

//BADD_813 replaced by BADD_830

//BADD_812 replaced by BADD_832

//BADD_811 replaced by BADD_831

//BADD_810 replaced by BADD_830

//KaratsubaCore_212 replaced by KaratsubaCore_230

//KaratsubaCore_211 replaced by KaratsubaCore_229

//KaratsubaCore_210 replaced by KaratsubaCore_228

//BADD_816 replaced by BADD_836

//BADD_815 replaced by BADD_835

//BADD_814 replaced by BADD_834

//KaratsubaCore_215 replaced by KaratsubaCore_233

//KaratsubaCore_214 replaced by KaratsubaCore_232

//KaratsubaCore_213 replaced by KaratsubaCore_231

//BADD_819 replaced by BADD_836

//BADD_818 replaced by BADD_835

//BADD_817 replaced by BADD_834

//KaratsubaCore_218 replaced by KaratsubaCore_233

//KaratsubaCore_217 replaced by KaratsubaCore_232

//KaratsubaCore_216 replaced by KaratsubaCore_231

//BADD_823 replaced by BADD_830

//BADD_822 replaced by BADD_832

//BADD_821 replaced by BADD_831

//BADD_820 replaced by BADD_830

//KaratsubaCore_221 replaced by KaratsubaCore_230

//KaratsubaCore_220 replaced by KaratsubaCore_229

//KaratsubaCore_219 replaced by KaratsubaCore_228

//BADD_826 replaced by BADD_836

//BADD_825 replaced by BADD_835

//BADD_824 replaced by BADD_834

//KaratsubaCore_224 replaced by KaratsubaCore_233

//KaratsubaCore_223 replaced by KaratsubaCore_232

//KaratsubaCore_222 replaced by KaratsubaCore_231

//BADD_829 replaced by BADD_836

//BADD_828 replaced by BADD_835

//BADD_827 replaced by BADD_834

//KaratsubaCore_227 replaced by KaratsubaCore_233

//KaratsubaCore_226 replaced by KaratsubaCore_232

//KaratsubaCore_225 replaced by KaratsubaCore_231

//BADD_833 replaced by BADD_830

module BADD_832 (
  input      [194:0]  io_a,
  input      [194:0]  io_b,
  input               io_c,
  output reg [195:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [48:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [48:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [3:0]    _zz__zz_io_s_12;
  wire       [3:0]    _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [3:0]    _zz_io_s_12;
  reg        [2:0]    _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,io_b[143 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {48'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,io_b[191 : 144]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {48'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[194 : 192]} + {1'b0,io_b[194 : 192]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {3'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[194 : 192] = _zz_io_s_13;
    io_s[195] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_13 <= _zz_io_s_12[2:0];
    _zz_io_s_14 <= _zz_io_s_12[3];
  end


endmodule

module BADD_831 (
  input      [194:0]  io_a,
  input      [194:0]  io_b,
  input               io_c,
  output reg [195:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [194:0]  _zz__zz_io_s_1;
  wire       [48:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [194:0]  _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_3_3;
  wire       [0:0]    _zz__zz_io_s_3_4;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [194:0]  _zz__zz_io_s_6_1;
  wire       [48:0]   _zz__zz_io_s_6_2;
  wire       [0:0]    _zz__zz_io_s_6_3;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [194:0]  _zz__zz_io_s_9_1;
  wire       [48:0]   _zz__zz_io_s_9_2;
  wire       [0:0]    _zz__zz_io_s_9_3;
  wire       [3:0]    _zz__zz_io_s_12;
  wire       [194:0]  _zz__zz_io_s_12_1;
  wire       [3:0]    _zz__zz_io_s_12_2;
  wire       [0:0]    _zz__zz_io_s_12_3;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [3:0]    _zz_io_s_12;
  reg        [2:0]    _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,_zz__zz_io_s_1[47 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {48'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_3_1 = ({1'b0,io_a[95 : 48]} + {1'b0,_zz__zz_io_s_3_2[95 : 48]});
  assign _zz__zz_io_s_3_2 = (~ io_b);
  assign _zz__zz_io_s_3_4 = _zz_io_s_2;
  assign _zz__zz_io_s_3_3 = {48'd0, _zz__zz_io_s_3_4};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,_zz__zz_io_s_6_1[143 : 96]});
  assign _zz__zz_io_s_6_1 = (~ io_b);
  assign _zz__zz_io_s_6_3 = _zz_io_s_5;
  assign _zz__zz_io_s_6_2 = {48'd0, _zz__zz_io_s_6_3};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,_zz__zz_io_s_9_1[191 : 144]});
  assign _zz__zz_io_s_9_1 = (~ io_b);
  assign _zz__zz_io_s_9_3 = _zz_io_s_8;
  assign _zz__zz_io_s_9_2 = {48'd0, _zz__zz_io_s_9_3};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[194 : 192]} + {1'b0,_zz__zz_io_s_12_1[194 : 192]});
  assign _zz__zz_io_s_12_1 = (~ io_b);
  assign _zz__zz_io_s_12_3 = _zz_io_s_11;
  assign _zz__zz_io_s_12_2 = {3'd0, _zz__zz_io_s_12_3};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[194 : 192] = _zz_io_s_13;
    io_s[195] = (! _zz_io_s_14);
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3_1 + _zz__zz_io_s_3_3);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_2);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_2);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_2);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_13 <= _zz_io_s_12[2:0];
    _zz_io_s_14 <= _zz_io_s_12[3];
  end


endmodule

module BADD_830 (
  input      [193:0]  io_a,
  input      [193:0]  io_b,
  input               io_c,
  output reg [194:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [48:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [48:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [2:0]    _zz__zz_io_s_12;
  wire       [2:0]    _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [2:0]    _zz_io_s_12;
  reg        [1:0]    _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,io_b[143 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {48'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,io_b[191 : 144]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {48'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[193 : 192]} + {1'b0,io_b[193 : 192]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {2'd0, _zz__zz_io_s_12_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[193 : 192] = _zz_io_s_13;
    io_s[194] = _zz_io_s_14;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_13 <= _zz_io_s_12[1:0];
    _zz_io_s_14 <= _zz_io_s_12[2];
  end


endmodule

module KaratsubaCore_230 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_a_1,
  input      [48:0]   io_b_0,
  input      [48:0]   io_b_1,
  output reg [193:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [98:0]   karatsuba_add2_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_b;
  wire       [97:0]   karatsuba_hasExtend_add4_io_a;
  wire       [97:0]   karatsuba_lsbMul_io_p;
  wire       [99:0]   karatsuba_midMul_io_p;
  wire       [97:0]   karatsuba_msbMul_io_p;
  wire       [98:0]   karatsuba_add1_io_s;
  wire       [99:0]   karatsuba_add2_io_s;
  wire       [99:0]   karatsuba_hasExtend_add3_io_s;
  wire       [98:0]   karatsuba_hasExtend_add4_io_s;
  wire       [51:0]   _zz_io_a;
  reg        [49:0]   _zz_io_a_0;
  reg        [49:0]   _zz_io_b_0;
  reg        [49:0]   _zz_io_b;
  reg        [97:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [97:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [97:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [97:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;

  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 48);
  KaratsubaCore_718 karatsuba_lsbMul (
    .io_a_0 (io_a_0[48:0]               ), //i
    .io_b_0 (io_b_0[48:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_715 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[49:0]           ), //i
    .io_b_0 (_zz_io_b_0[49:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_718 karatsuba_msbMul (
    .io_a_0 (io_a_1[48:0]               ), //i
    .io_b_0 (io_b_1[48:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1406 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[97:0]), //i
    .io_b   (karatsuba_msbMul_io_p[97:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[98:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1407 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[98:0]), //i
    .io_b   (karatsuba_add1_io_s[98:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[99:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_1408 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[98:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[98:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[99:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  BADD_1406 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[97:0]                 ), //i
    .io_b   (karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4[97:0]), //i
    .io_c   (1'b0                                                ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[98:0]                 ), //o
    .clk    (clk                                                 ), //i
    .resetn (resetn                                              )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[98:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[98:0];
  assign karatsuba_hasExtend_add3_io_b = {49'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {46'd0, _zz_io_a};
  always @(*) begin
    io_p[47 : 0] = _zz_io_p_2;
    io_p[95 : 48] = _zz_io_p_3;
    io_p[193 : 96] = karatsuba_hasExtend_add4_io_s[97:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_1});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_1});
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= karatsuba_hasExtend_add3_io_s[47:0];
  end


endmodule

module KaratsubaCore_229 (
  input      [49:0]   io_a_0,
  input      [49:0]   io_a_1,
  input      [49:0]   io_b_0,
  input      [49:0]   io_b_1,
  output reg [195:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [100:0]  karatsuba_add2_io_a;
  wire       [100:0]  karatsuba_hasExtend_add3_io_a;
  wire       [100:0]  karatsuba_hasExtend_add3_io_b;
  wire       [99:0]   karatsuba_hasExtend_add4_io_a;
  wire       [99:0]   karatsuba_lsbMul_io_p;
  wire       [101:0]  karatsuba_midMul_io_p;
  wire       [99:0]   karatsuba_msbMul_io_p;
  wire       [100:0]  karatsuba_add1_io_s;
  wire       [101:0]  karatsuba_add2_io_s;
  wire       [101:0]  karatsuba_hasExtend_add3_io_s;
  wire       [100:0]  karatsuba_hasExtend_add4_io_s;
  wire       [53:0]   _zz_io_a;
  reg        [50:0]   _zz_io_a_0;
  reg        [50:0]   _zz_io_b_0;
  reg        [51:0]   _zz_io_b;
  reg        [99:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
  reg        [99:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
  reg        [99:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
  reg        [99:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_4;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;

  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 48);
  KaratsubaCore_715 karatsuba_lsbMul (
    .io_a_0 (io_a_0[49:0]               ), //i
    .io_b_0 (io_b_0[49:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_706 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[50:0]            ), //i
    .io_b_0 (_zz_io_b_0[50:0]            ), //i
    .io_p   (karatsuba_midMul_io_p[101:0]), //o
    .clk    (clk                         ), //i
    .resetn (resetn                      )  //i
  );
  KaratsubaCore_715 karatsuba_msbMul (
    .io_a_0 (io_a_1[49:0]               ), //i
    .io_b_0 (io_b_1[49:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1395 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[99:0]), //i
    .io_b   (karatsuba_msbMul_io_p[99:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[100:0] ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1396 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[100:0]), //i
    .io_b   (karatsuba_add1_io_s[100:0]), //i
    .io_c   (1'b1                      ), //i
    .io_s   (karatsuba_add2_io_s[101:0]), //o
    .clk    (clk                       ), //i
    .resetn (resetn                    )  //i
  );
  BADD_1397 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[100:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[100:0]), //i
    .io_c   (1'b0                                ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[101:0]), //o
    .clk    (clk                                 ), //i
    .resetn (resetn                              )  //i
  );
  BADD_1395 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[99:0]                 ), //i
    .io_b   (karatsuba_midMul_karatsuba_msbMul_io_p_delay_4[99:0]), //i
    .io_c   (1'b0                                                ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[100:0]                ), //o
    .clk    (clk                                                 ), //i
    .resetn (resetn                                              )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[100:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[100:0];
  assign karatsuba_hasExtend_add3_io_b = {49'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {46'd0, _zz_io_a};
  always @(*) begin
    io_p[47 : 0] = _zz_io_p_2;
    io_p[95 : 48] = _zz_io_p_3;
    io_p[195 : 96] = karatsuba_hasExtend_add4_io_s[99:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_1});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_1});
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= karatsuba_hasExtend_add3_io_s[47:0];
  end


endmodule

module KaratsubaCore_228 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_a_1,
  input      [48:0]   io_b_0,
  input      [48:0]   io_b_1,
  output reg [193:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [98:0]   karatsuba_add2_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_b;
  wire       [97:0]   karatsuba_hasExtend_add4_io_a;
  wire       [97:0]   karatsuba_lsbMul_io_p;
  wire       [99:0]   karatsuba_midMul_io_p;
  wire       [97:0]   karatsuba_msbMul_io_p;
  wire       [98:0]   karatsuba_add1_io_s;
  wire       [99:0]   karatsuba_add2_io_s;
  wire       [99:0]   karatsuba_hasExtend_add3_io_s;
  wire       [98:0]   karatsuba_hasExtend_add4_io_s;
  wire       [51:0]   _zz_io_a;
  reg        [49:0]   _zz_io_a_0;
  reg        [49:0]   _zz_io_b_0;
  reg        [49:0]   _zz_io_b;
  reg        [97:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [97:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [97:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [97:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;

  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 48);
  KaratsubaCore_718 karatsuba_lsbMul (
    .io_a_0 (io_a_0[48:0]               ), //i
    .io_b_0 (io_b_0[48:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_715 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[49:0]           ), //i
    .io_b_0 (_zz_io_b_0[49:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_718 karatsuba_msbMul (
    .io_a_0 (io_a_1[48:0]               ), //i
    .io_b_0 (io_b_1[48:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1406 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[97:0]), //i
    .io_b   (karatsuba_msbMul_io_p[97:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[98:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1407 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[98:0]), //i
    .io_b   (karatsuba_add1_io_s[98:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[99:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_1408 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[98:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[98:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[99:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  BADD_1406 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[97:0]                 ), //i
    .io_b   (karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4[97:0]), //i
    .io_c   (1'b0                                                ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[98:0]                 ), //o
    .clk    (clk                                                 ), //i
    .resetn (resetn                                              )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[98:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[98:0];
  assign karatsuba_hasExtend_add3_io_b = {49'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {46'd0, _zz_io_a};
  always @(*) begin
    io_p[47 : 0] = _zz_io_p_2;
    io_p[95 : 48] = _zz_io_p_3;
    io_p[193 : 96] = karatsuba_hasExtend_add4_io_s[97:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_1});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_1});
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= karatsuba_hasExtend_add3_io_s[47:0];
  end


endmodule

module BADD_836 (
  input      [287:0]  io_a,
  input      [287:0]  io_b,
  input               io_c,
  output reg [288:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [48:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [48:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [48:0]   _zz__zz_io_s_12;
  wire       [48:0]   _zz__zz_io_s_12_1;
  wire       [0:0]    _zz__zz_io_s_12_2;
  wire       [48:0]   _zz__zz_io_s_15;
  wire       [48:0]   _zz__zz_io_s_15_1;
  wire       [0:0]    _zz__zz_io_s_15_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [48:0]   _zz_io_s_12;
  reg        [47:0]   _zz_io_s_13;
  reg                 _zz_io_s_14;
  wire       [48:0]   _zz_io_s_15;
  reg        [47:0]   _zz_io_s_16;
  reg                 _zz_io_s_17;
  reg                 _zz_io_s_18;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,io_b[143 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {48'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,io_b[191 : 144]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {48'd0, _zz__zz_io_s_9_2};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[239 : 192]} + {1'b0,io_b[239 : 192]});
  assign _zz__zz_io_s_12_2 = _zz_io_s_11;
  assign _zz__zz_io_s_12_1 = {48'd0, _zz__zz_io_s_12_2};
  assign _zz__zz_io_s_15 = ({1'b0,io_a[287 : 240]} + {1'b0,io_b[287 : 240]});
  assign _zz__zz_io_s_15_2 = _zz_io_s_14;
  assign _zz__zz_io_s_15_1 = {48'd0, _zz__zz_io_s_15_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[239 : 192] = _zz_io_s_13;
    io_s[287 : 240] = _zz_io_s_16;
    io_s[288] = _zz_io_s_18;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_1);
  assign _zz_io_s_15 = (_zz__zz_io_s_15 + _zz__zz_io_s_15_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_13 <= _zz_io_s_12[47:0];
    _zz_io_s_14 <= _zz_io_s_12[48];
    _zz_io_s_16 <= _zz_io_s_15[47:0];
    _zz_io_s_17 <= _zz_io_s_15[48];
    _zz_io_s_18 <= _zz_io_s_17;
  end


endmodule

module BADD_835 (
  input      [192:0]  io_a,
  input      [192:0]  io_b,
  input               io_c,
  output reg [193:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [192:0]  _zz__zz_io_s_1;
  wire       [48:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [192:0]  _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_3_3;
  wire       [0:0]    _zz__zz_io_s_3_4;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [192:0]  _zz__zz_io_s_6_1;
  wire       [48:0]   _zz__zz_io_s_6_2;
  wire       [0:0]    _zz__zz_io_s_6_3;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [192:0]  _zz__zz_io_s_9_1;
  wire       [48:0]   _zz__zz_io_s_9_2;
  wire       [0:0]    _zz__zz_io_s_9_3;
  wire       [1:0]    _zz__zz_io_s_12;
  wire       [192:0]  _zz__zz_io_s_12_1;
  wire       [1:0]    _zz__zz_io_s_12_2;
  wire       [0:0]    _zz__zz_io_s_12_3;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  wire       [1:0]    _zz_io_s_12;
  reg        [0:0]    _zz_io_s_13;
  reg                 _zz_io_s_14;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,_zz__zz_io_s_1[47 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {48'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_3_1 = ({1'b0,io_a[95 : 48]} + {1'b0,_zz__zz_io_s_3_2[95 : 48]});
  assign _zz__zz_io_s_3_2 = (~ io_b);
  assign _zz__zz_io_s_3_4 = _zz_io_s_2;
  assign _zz__zz_io_s_3_3 = {48'd0, _zz__zz_io_s_3_4};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,_zz__zz_io_s_6_1[143 : 96]});
  assign _zz__zz_io_s_6_1 = (~ io_b);
  assign _zz__zz_io_s_6_3 = _zz_io_s_5;
  assign _zz__zz_io_s_6_2 = {48'd0, _zz__zz_io_s_6_3};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,_zz__zz_io_s_9_1[191 : 144]});
  assign _zz__zz_io_s_9_1 = (~ io_b);
  assign _zz__zz_io_s_9_3 = _zz_io_s_8;
  assign _zz__zz_io_s_9_2 = {48'd0, _zz__zz_io_s_9_3};
  assign _zz__zz_io_s_12 = ({1'b0,io_a[192 : 192]} + {1'b0,_zz__zz_io_s_12_1[192 : 192]});
  assign _zz__zz_io_s_12_1 = (~ io_b);
  assign _zz__zz_io_s_12_3 = _zz_io_s_11;
  assign _zz__zz_io_s_12_2 = {1'd0, _zz__zz_io_s_12_3};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[192 : 192] = _zz_io_s_13;
    io_s[193] = (! _zz_io_s_14);
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3_1 + _zz__zz_io_s_3_3);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_2);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_2);
  assign _zz_io_s_12 = (_zz__zz_io_s_12 + _zz__zz_io_s_12_2);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_13 <= _zz_io_s_12[0:0];
    _zz_io_s_14 <= _zz_io_s_12[1];
  end


endmodule

module BADD_834 (
  input      [191:0]  io_a,
  input      [191:0]  io_b,
  input               io_c,
  output reg [192:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [48:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz__zz_io_s_9;
  wire       [48:0]   _zz__zz_io_s_9_1;
  wire       [0:0]    _zz__zz_io_s_9_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  wire       [48:0]   _zz_io_s_9;
  reg        [47:0]   _zz_io_s_10;
  reg                 _zz_io_s_11;
  reg                 _zz_io_s_12;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,io_b[143 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {48'd0, _zz__zz_io_s_6_2};
  assign _zz__zz_io_s_9 = ({1'b0,io_a[191 : 144]} + {1'b0,io_b[191 : 144]});
  assign _zz__zz_io_s_9_2 = _zz_io_s_8;
  assign _zz__zz_io_s_9_1 = {48'd0, _zz__zz_io_s_9_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[191 : 144] = _zz_io_s_10;
    io_s[192] = _zz_io_s_12;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  assign _zz_io_s_9 = (_zz__zz_io_s_9 + _zz__zz_io_s_9_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_10 <= _zz_io_s_9[47:0];
    _zz_io_s_11 <= _zz_io_s_9[48];
    _zz_io_s_12 <= _zz_io_s_11;
  end


endmodule

module KaratsubaCore_233 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  output reg [191:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [96:0]   karatsuba_add2_io_a;
  wire       [143:0]  karatsuba_noExtend_add3_io_a;
  reg        [143:0]  karatsuba_noExtend_add3_io_b;
  wire       [95:0]   karatsuba_lsbMul_io_p;
  wire       [97:0]   karatsuba_midMul_io_p;
  wire       [95:0]   karatsuba_msbMul_io_p;
  wire       [96:0]   karatsuba_add1_io_s;
  wire       [97:0]   karatsuba_add2_io_s;
  wire       [144:0]  karatsuba_noExtend_add3_io_s;
  wire       [96:0]   _zz_io_a;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_b_0;
  reg        [47:0]   _zz_io_b;
  reg        [95:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [95:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [95:0]   karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;

  assign _zz_io_a = karatsuba_add2_io_s[96:0];
  KaratsubaCore_717 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]               ), //i
    .io_b_0 (io_b_0[47:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[95:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_718 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]           ), //i
    .io_b_0 (_zz_io_b_0[48:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_717 karatsuba_msbMul (
    .io_a_0 (io_a_1[47:0]               ), //i
    .io_b_0 (io_b_1[47:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[95:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1410 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[95:0]), //i
    .io_b   (karatsuba_msbMul_io_p[95:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[96:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1411 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[96:0]), //i
    .io_b   (karatsuba_add1_io_s[96:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[97:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_1412 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[143:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[143:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[144:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[96:0];
  assign karatsuba_noExtend_add3_io_a = {47'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[47 : 0] = _zz_io_b;
    karatsuba_noExtend_add3_io_b[143 : 48] = karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3;
  end

  always @(*) begin
    io_p[47 : 0] = _zz_io_p_1;
    io_p[191 : 48] = karatsuba_noExtend_add3_io_s[143:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_1});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_1});
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_msbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_msbMul_karatsuba_msbMul_io_p_delay_2;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
  end


endmodule

module KaratsubaCore_232 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_a_1,
  input      [48:0]   io_b_0,
  input      [48:0]   io_b_1,
  output reg [193:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [98:0]   karatsuba_add2_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_a;
  wire       [98:0]   karatsuba_hasExtend_add3_io_b;
  wire       [97:0]   karatsuba_hasExtend_add4_io_a;
  wire       [97:0]   karatsuba_lsbMul_io_p;
  wire       [99:0]   karatsuba_midMul_io_p;
  wire       [97:0]   karatsuba_msbMul_io_p;
  wire       [98:0]   karatsuba_add1_io_s;
  wire       [99:0]   karatsuba_add2_io_s;
  wire       [99:0]   karatsuba_hasExtend_add3_io_s;
  wire       [98:0]   karatsuba_hasExtend_add4_io_s;
  wire       [51:0]   _zz_io_a;
  reg        [49:0]   _zz_io_a_0;
  reg        [49:0]   _zz_io_b_0;
  reg        [49:0]   _zz_io_b;
  reg        [97:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
  reg        [97:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
  reg        [97:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
  reg        [97:0]   karatsuba_midMul_karatsuba_msbMul_io_p_delay_4;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;
  reg        [47:0]   _zz_io_p_2;
  reg        [47:0]   _zz_io_p_3;

  assign _zz_io_a = (karatsuba_hasExtend_add3_io_s >>> 48);
  KaratsubaCore_718 karatsuba_lsbMul (
    .io_a_0 (io_a_0[48:0]               ), //i
    .io_b_0 (io_b_0[48:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_715 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[49:0]           ), //i
    .io_b_0 (_zz_io_b_0[49:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[99:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_718 karatsuba_msbMul (
    .io_a_0 (io_a_1[48:0]               ), //i
    .io_b_0 (io_b_1[48:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1406 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[97:0]), //i
    .io_b   (karatsuba_msbMul_io_p[97:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[98:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1407 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[98:0]), //i
    .io_b   (karatsuba_add1_io_s[98:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[99:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_1408 karatsuba_hasExtend_add3 (
    .io_a   (karatsuba_hasExtend_add3_io_a[98:0]), //i
    .io_b   (karatsuba_hasExtend_add3_io_b[98:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_hasExtend_add3_io_s[99:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  BADD_1406 karatsuba_hasExtend_add4 (
    .io_a   (karatsuba_hasExtend_add4_io_a[97:0]                 ), //i
    .io_b   (karatsuba_midMul_karatsuba_msbMul_io_p_delay_4[97:0]), //i
    .io_c   (1'b0                                                ), //i
    .io_s   (karatsuba_hasExtend_add4_io_s[98:0]                 ), //o
    .clk    (clk                                                 ), //i
    .resetn (resetn                                              )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[98:0];
  assign karatsuba_hasExtend_add3_io_a = karatsuba_add2_io_s[98:0];
  assign karatsuba_hasExtend_add3_io_b = {49'd0, _zz_io_b};
  assign karatsuba_hasExtend_add4_io_a = {46'd0, _zz_io_a};
  always @(*) begin
    io_p[47 : 0] = _zz_io_p_2;
    io_p[95 : 48] = _zz_io_p_3;
    io_p[193 : 96] = karatsuba_hasExtend_add4_io_s[97:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_1});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_1});
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_2;
    karatsuba_midMul_karatsuba_msbMul_io_p_delay_4 <= karatsuba_midMul_karatsuba_msbMul_io_p_delay_3;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= karatsuba_hasExtend_add3_io_s[47:0];
  end


endmodule

module KaratsubaCore_231 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_a_1,
  input      [47:0]   io_b_0,
  input      [47:0]   io_b_1,
  output reg [191:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [96:0]   karatsuba_add2_io_a;
  wire       [143:0]  karatsuba_noExtend_add3_io_a;
  reg        [143:0]  karatsuba_noExtend_add3_io_b;
  wire       [95:0]   karatsuba_lsbMul_io_p;
  wire       [97:0]   karatsuba_midMul_io_p;
  wire       [95:0]   karatsuba_msbMul_io_p;
  wire       [96:0]   karatsuba_add1_io_s;
  wire       [97:0]   karatsuba_add2_io_s;
  wire       [144:0]  karatsuba_noExtend_add3_io_s;
  wire       [96:0]   _zz_io_a;
  reg        [48:0]   _zz_io_a_0;
  reg        [48:0]   _zz_io_b_0;
  reg        [47:0]   _zz_io_b;
  reg        [95:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
  reg        [95:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
  reg        [95:0]   karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
  reg        [47:0]   _zz_io_p;
  reg        [47:0]   _zz_io_p_1;

  assign _zz_io_a = karatsuba_add2_io_s[96:0];
  KaratsubaCore_717 karatsuba_lsbMul (
    .io_a_0 (io_a_0[47:0]               ), //i
    .io_b_0 (io_b_0[47:0]               ), //i
    .io_p   (karatsuba_lsbMul_io_p[95:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_718 karatsuba_midMul (
    .io_a_0 (_zz_io_a_0[48:0]           ), //i
    .io_b_0 (_zz_io_b_0[48:0]           ), //i
    .io_p   (karatsuba_midMul_io_p[97:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  KaratsubaCore_717 karatsuba_msbMul (
    .io_a_0 (io_a_1[47:0]               ), //i
    .io_b_0 (io_b_1[47:0]               ), //i
    .io_p   (karatsuba_msbMul_io_p[95:0]), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1410 karatsuba_add1 (
    .io_a   (karatsuba_lsbMul_io_p[95:0]), //i
    .io_b   (karatsuba_msbMul_io_p[95:0]), //i
    .io_c   (1'b0                       ), //i
    .io_s   (karatsuba_add1_io_s[96:0]  ), //o
    .clk    (clk                        ), //i
    .resetn (resetn                     )  //i
  );
  BADD_1411 karatsuba_add2 (
    .io_a   (karatsuba_add2_io_a[96:0]), //i
    .io_b   (karatsuba_add1_io_s[96:0]), //i
    .io_c   (1'b1                     ), //i
    .io_s   (karatsuba_add2_io_s[97:0]), //o
    .clk    (clk                      ), //i
    .resetn (resetn                   )  //i
  );
  BADD_1412 karatsuba_noExtend_add3 (
    .io_a   (karatsuba_noExtend_add3_io_a[143:0]), //i
    .io_b   (karatsuba_noExtend_add3_io_b[143:0]), //i
    .io_c   (1'b0                               ), //i
    .io_s   (karatsuba_noExtend_add3_io_s[144:0]), //o
    .clk    (clk                                ), //i
    .resetn (resetn                             )  //i
  );
  assign karatsuba_add2_io_a = karatsuba_midMul_io_p[96:0];
  assign karatsuba_noExtend_add3_io_a = {47'd0, _zz_io_a};
  always @(*) begin
    karatsuba_noExtend_add3_io_b[47 : 0] = _zz_io_b;
    karatsuba_noExtend_add3_io_b[143 : 48] = karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3;
  end

  always @(*) begin
    io_p[47 : 0] = _zz_io_p_1;
    io_p[191 : 48] = karatsuba_noExtend_add3_io_s[143:0];
  end

  always @(posedge clk) begin
    _zz_io_a_0 <= ({1'b0,io_a_0} + {1'b0,io_a_1});
    _zz_io_b_0 <= ({1'b0,io_b_0} + {1'b0,io_b_1});
    _zz_io_b <= (karatsuba_lsbMul_io_p >>> 48);
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1 <= karatsuba_msbMul_io_p;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_1;
    karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_3 <= karatsuba_lsbMul_karatsuba_msbMul_io_p_delay_2;
    _zz_io_p <= karatsuba_lsbMul_io_p[47 : 0];
    _zz_io_p_1 <= _zz_io_p;
  end


endmodule

//BADD_839 replaced by BADD_1412

//BADD_838 replaced by BADD_1411

//BADD_837 replaced by BADD_1410

//KaratsubaCore_236 replaced by KaratsubaCore_717

//KaratsubaCore_235 replaced by KaratsubaCore_718

//KaratsubaCore_234 replaced by KaratsubaCore_717

//BADD_843 replaced by BADD_1406

//BADD_842 replaced by BADD_1408

//BADD_841 replaced by BADD_1407

//BADD_840 replaced by BADD_1406

//KaratsubaCore_239 replaced by KaratsubaCore_718

//KaratsubaCore_238 replaced by KaratsubaCore_715

//KaratsubaCore_237 replaced by KaratsubaCore_718

//BADD_846 replaced by BADD_1412

//BADD_845 replaced by BADD_1411

//BADD_844 replaced by BADD_1410

//KaratsubaCore_242 replaced by KaratsubaCore_717

//KaratsubaCore_241 replaced by KaratsubaCore_718

//KaratsubaCore_240 replaced by KaratsubaCore_717

//BADD_850 replaced by BADD_1406

//BADD_849 replaced by BADD_1408

//BADD_848 replaced by BADD_1407

//BADD_847 replaced by BADD_1406

//KaratsubaCore_245 replaced by KaratsubaCore_718

//KaratsubaCore_244 replaced by KaratsubaCore_715

//KaratsubaCore_243 replaced by KaratsubaCore_718

//BADD_854 replaced by BADD_1395

//BADD_853 replaced by BADD_1397

//BADD_852 replaced by BADD_1396

//BADD_851 replaced by BADD_1395

//KaratsubaCore_248 replaced by KaratsubaCore_715

//KaratsubaCore_247 replaced by KaratsubaCore_706

//KaratsubaCore_246 replaced by KaratsubaCore_715

//BADD_858 replaced by BADD_1406

//BADD_857 replaced by BADD_1408

//BADD_856 replaced by BADD_1407

//BADD_855 replaced by BADD_1406

//KaratsubaCore_251 replaced by KaratsubaCore_718

//KaratsubaCore_250 replaced by KaratsubaCore_715

//KaratsubaCore_249 replaced by KaratsubaCore_718

//BADD_861 replaced by BADD_1412

//BADD_860 replaced by BADD_1411

//BADD_859 replaced by BADD_1410

//KaratsubaCore_254 replaced by KaratsubaCore_717

//KaratsubaCore_253 replaced by KaratsubaCore_718

//KaratsubaCore_252 replaced by KaratsubaCore_717

//BADD_865 replaced by BADD_1406

//BADD_864 replaced by BADD_1408

//BADD_863 replaced by BADD_1407

//BADD_862 replaced by BADD_1406

//KaratsubaCore_257 replaced by KaratsubaCore_718

//KaratsubaCore_256 replaced by KaratsubaCore_715

//KaratsubaCore_255 replaced by KaratsubaCore_718

//BADD_868 replaced by BADD_1412

//BADD_867 replaced by BADD_1411

//BADD_866 replaced by BADD_1410

//KaratsubaCore_260 replaced by KaratsubaCore_717

//KaratsubaCore_259 replaced by KaratsubaCore_718

//KaratsubaCore_258 replaced by KaratsubaCore_717

//BADD_871 replaced by BADD_1412

//BADD_870 replaced by BADD_1411

//BADD_869 replaced by BADD_1410

//KaratsubaCore_263 replaced by KaratsubaCore_717

//KaratsubaCore_262 replaced by KaratsubaCore_718

//KaratsubaCore_261 replaced by KaratsubaCore_717

//BADD_875 replaced by BADD_1406

//BADD_874 replaced by BADD_1408

//BADD_873 replaced by BADD_1407

//BADD_872 replaced by BADD_1406

//KaratsubaCore_266 replaced by KaratsubaCore_718

//KaratsubaCore_265 replaced by KaratsubaCore_715

//KaratsubaCore_264 replaced by KaratsubaCore_718

//BADD_878 replaced by BADD_1412

//BADD_877 replaced by BADD_1411

//BADD_876 replaced by BADD_1410

//KaratsubaCore_269 replaced by KaratsubaCore_717

//KaratsubaCore_268 replaced by KaratsubaCore_718

//KaratsubaCore_267 replaced by KaratsubaCore_717

//BADD_882 replaced by BADD_1406

//BADD_881 replaced by BADD_1408

//BADD_880 replaced by BADD_1407

//BADD_879 replaced by BADD_1406

//KaratsubaCore_272 replaced by KaratsubaCore_718

//KaratsubaCore_271 replaced by KaratsubaCore_715

//KaratsubaCore_270 replaced by KaratsubaCore_718

//BADD_886 replaced by BADD_1395

//BADD_885 replaced by BADD_1397

//BADD_884 replaced by BADD_1396

//BADD_883 replaced by BADD_1395

//KaratsubaCore_275 replaced by KaratsubaCore_715

//KaratsubaCore_274 replaced by KaratsubaCore_706

//KaratsubaCore_273 replaced by KaratsubaCore_715

//BADD_890 replaced by BADD_1406

//BADD_889 replaced by BADD_1408

//BADD_888 replaced by BADD_1407

//BADD_887 replaced by BADD_1406

//KaratsubaCore_278 replaced by KaratsubaCore_718

//KaratsubaCore_277 replaced by KaratsubaCore_715

//KaratsubaCore_276 replaced by KaratsubaCore_718

//BADD_893 replaced by BADD_1412

//BADD_892 replaced by BADD_1411

//BADD_891 replaced by BADD_1410

//KaratsubaCore_281 replaced by KaratsubaCore_717

//KaratsubaCore_280 replaced by KaratsubaCore_718

//KaratsubaCore_279 replaced by KaratsubaCore_717

//BADD_897 replaced by BADD_1406

//BADD_896 replaced by BADD_1408

//BADD_895 replaced by BADD_1407

//BADD_894 replaced by BADD_1406

//KaratsubaCore_284 replaced by KaratsubaCore_718

//KaratsubaCore_283 replaced by KaratsubaCore_715

//KaratsubaCore_282 replaced by KaratsubaCore_718

//BADD_900 replaced by BADD_1412

//BADD_899 replaced by BADD_1411

//BADD_898 replaced by BADD_1410

//KaratsubaCore_287 replaced by KaratsubaCore_717

//KaratsubaCore_286 replaced by KaratsubaCore_718

//KaratsubaCore_285 replaced by KaratsubaCore_717

//BADD_903 replaced by BADD_1412

//BADD_902 replaced by BADD_1411

//BADD_901 replaced by BADD_1410

//KaratsubaCore_290 replaced by KaratsubaCore_717

//KaratsubaCore_289 replaced by KaratsubaCore_718

//KaratsubaCore_288 replaced by KaratsubaCore_717

//BADD_907 replaced by BADD_1406

//BADD_906 replaced by BADD_1408

//BADD_905 replaced by BADD_1407

//BADD_904 replaced by BADD_1406

//KaratsubaCore_293 replaced by KaratsubaCore_718

//KaratsubaCore_292 replaced by KaratsubaCore_715

//KaratsubaCore_291 replaced by KaratsubaCore_718

//BADD_910 replaced by BADD_1412

//BADD_909 replaced by BADD_1411

//BADD_908 replaced by BADD_1410

//KaratsubaCore_296 replaced by KaratsubaCore_717

//KaratsubaCore_295 replaced by KaratsubaCore_718

//KaratsubaCore_294 replaced by KaratsubaCore_717

//BADD_914 replaced by BADD_1406

//BADD_913 replaced by BADD_1408

//BADD_912 replaced by BADD_1407

//BADD_911 replaced by BADD_1406

//KaratsubaCore_299 replaced by KaratsubaCore_718

//KaratsubaCore_298 replaced by KaratsubaCore_715

//KaratsubaCore_297 replaced by KaratsubaCore_718

//BADD_918 replaced by BADD_1395

//BADD_917 replaced by BADD_1397

//BADD_916 replaced by BADD_1396

//BADD_915 replaced by BADD_1395

//KaratsubaCore_302 replaced by KaratsubaCore_715

//KaratsubaCore_301 replaced by KaratsubaCore_706

//KaratsubaCore_300 replaced by KaratsubaCore_715

//BADD_922 replaced by BADD_1406

//BADD_921 replaced by BADD_1408

//BADD_920 replaced by BADD_1407

//BADD_919 replaced by BADD_1406

//KaratsubaCore_305 replaced by KaratsubaCore_718

//KaratsubaCore_304 replaced by KaratsubaCore_715

//KaratsubaCore_303 replaced by KaratsubaCore_718

//BADD_925 replaced by BADD_1412

//BADD_924 replaced by BADD_1411

//BADD_923 replaced by BADD_1410

//KaratsubaCore_308 replaced by KaratsubaCore_717

//KaratsubaCore_307 replaced by KaratsubaCore_718

//KaratsubaCore_306 replaced by KaratsubaCore_717

//BADD_929 replaced by BADD_1406

//BADD_928 replaced by BADD_1408

//BADD_927 replaced by BADD_1407

//BADD_926 replaced by BADD_1406

//KaratsubaCore_311 replaced by KaratsubaCore_718

//KaratsubaCore_310 replaced by KaratsubaCore_715

//KaratsubaCore_309 replaced by KaratsubaCore_718

//BADD_932 replaced by BADD_1412

//BADD_931 replaced by BADD_1411

//BADD_930 replaced by BADD_1410

//KaratsubaCore_314 replaced by KaratsubaCore_717

//KaratsubaCore_313 replaced by KaratsubaCore_718

//KaratsubaCore_312 replaced by KaratsubaCore_717

//BADD_935 replaced by BADD_1412

//BADD_934 replaced by BADD_1411

//BADD_933 replaced by BADD_1410

//KaratsubaCore_317 replaced by KaratsubaCore_717

//KaratsubaCore_316 replaced by KaratsubaCore_718

//KaratsubaCore_315 replaced by KaratsubaCore_717

//BADD_939 replaced by BADD_1406

//BADD_938 replaced by BADD_1408

//BADD_937 replaced by BADD_1407

//BADD_936 replaced by BADD_1406

//KaratsubaCore_320 replaced by KaratsubaCore_718

//KaratsubaCore_319 replaced by KaratsubaCore_715

//KaratsubaCore_318 replaced by KaratsubaCore_718

//BADD_942 replaced by BADD_1412

//BADD_941 replaced by BADD_1411

//BADD_940 replaced by BADD_1410

//KaratsubaCore_323 replaced by KaratsubaCore_717

//KaratsubaCore_322 replaced by KaratsubaCore_718

//KaratsubaCore_321 replaced by KaratsubaCore_717

//BADD_946 replaced by BADD_1406

//BADD_945 replaced by BADD_1408

//BADD_944 replaced by BADD_1407

//BADD_943 replaced by BADD_1406

//KaratsubaCore_326 replaced by KaratsubaCore_718

//KaratsubaCore_325 replaced by KaratsubaCore_715

//KaratsubaCore_324 replaced by KaratsubaCore_718

//BADD_950 replaced by BADD_1395

//BADD_949 replaced by BADD_1397

//BADD_948 replaced by BADD_1396

//BADD_947 replaced by BADD_1395

//KaratsubaCore_329 replaced by KaratsubaCore_715

//KaratsubaCore_328 replaced by KaratsubaCore_706

//KaratsubaCore_327 replaced by KaratsubaCore_715

//BADD_954 replaced by BADD_1406

//BADD_953 replaced by BADD_1408

//BADD_952 replaced by BADD_1407

//BADD_951 replaced by BADD_1406

//KaratsubaCore_332 replaced by KaratsubaCore_718

//KaratsubaCore_331 replaced by KaratsubaCore_715

//KaratsubaCore_330 replaced by KaratsubaCore_718

//BADD_957 replaced by BADD_1412

//BADD_956 replaced by BADD_1411

//BADD_955 replaced by BADD_1410

//KaratsubaCore_335 replaced by KaratsubaCore_717

//KaratsubaCore_334 replaced by KaratsubaCore_718

//KaratsubaCore_333 replaced by KaratsubaCore_717

//BADD_961 replaced by BADD_1406

//BADD_960 replaced by BADD_1408

//BADD_959 replaced by BADD_1407

//BADD_958 replaced by BADD_1406

//KaratsubaCore_338 replaced by KaratsubaCore_718

//KaratsubaCore_337 replaced by KaratsubaCore_715

//KaratsubaCore_336 replaced by KaratsubaCore_718

//BADD_964 replaced by BADD_1412

//BADD_963 replaced by BADD_1411

//BADD_962 replaced by BADD_1410

//KaratsubaCore_341 replaced by KaratsubaCore_717

//KaratsubaCore_340 replaced by KaratsubaCore_718

//KaratsubaCore_339 replaced by KaratsubaCore_717

//BADD_967 replaced by BADD_1412

//BADD_966 replaced by BADD_1411

//BADD_965 replaced by BADD_1410

//KaratsubaCore_344 replaced by KaratsubaCore_717

//KaratsubaCore_343 replaced by KaratsubaCore_718

//KaratsubaCore_342 replaced by KaratsubaCore_717

//BADD_971 replaced by BADD_1406

//BADD_970 replaced by BADD_1408

//BADD_969 replaced by BADD_1407

//BADD_968 replaced by BADD_1406

//KaratsubaCore_347 replaced by KaratsubaCore_718

//KaratsubaCore_346 replaced by KaratsubaCore_715

//KaratsubaCore_345 replaced by KaratsubaCore_718

//BADD_974 replaced by BADD_1412

//BADD_973 replaced by BADD_1411

//BADD_972 replaced by BADD_1410

//KaratsubaCore_350 replaced by KaratsubaCore_717

//KaratsubaCore_349 replaced by KaratsubaCore_718

//KaratsubaCore_348 replaced by KaratsubaCore_717

//BADD_978 replaced by BADD_1406

//BADD_977 replaced by BADD_1408

//BADD_976 replaced by BADD_1407

//BADD_975 replaced by BADD_1406

//KaratsubaCore_353 replaced by KaratsubaCore_718

//KaratsubaCore_352 replaced by KaratsubaCore_715

//KaratsubaCore_351 replaced by KaratsubaCore_718

//BADD_982 replaced by BADD_1395

//BADD_981 replaced by BADD_1397

//BADD_980 replaced by BADD_1396

//BADD_979 replaced by BADD_1395

//KaratsubaCore_356 replaced by KaratsubaCore_715

//KaratsubaCore_355 replaced by KaratsubaCore_706

//KaratsubaCore_354 replaced by KaratsubaCore_715

//BADD_986 replaced by BADD_1406

//BADD_985 replaced by BADD_1408

//BADD_984 replaced by BADD_1407

//BADD_983 replaced by BADD_1406

//KaratsubaCore_359 replaced by KaratsubaCore_718

//KaratsubaCore_358 replaced by KaratsubaCore_715

//KaratsubaCore_357 replaced by KaratsubaCore_718

//BADD_989 replaced by BADD_1412

//BADD_988 replaced by BADD_1411

//BADD_987 replaced by BADD_1410

//KaratsubaCore_362 replaced by KaratsubaCore_717

//KaratsubaCore_361 replaced by KaratsubaCore_718

//KaratsubaCore_360 replaced by KaratsubaCore_717

//BADD_993 replaced by BADD_1406

//BADD_992 replaced by BADD_1408

//BADD_991 replaced by BADD_1407

//BADD_990 replaced by BADD_1406

//KaratsubaCore_365 replaced by KaratsubaCore_718

//KaratsubaCore_364 replaced by KaratsubaCore_715

//KaratsubaCore_363 replaced by KaratsubaCore_718

//BADD_996 replaced by BADD_1412

//BADD_995 replaced by BADD_1411

//BADD_994 replaced by BADD_1410

//KaratsubaCore_368 replaced by KaratsubaCore_717

//KaratsubaCore_367 replaced by KaratsubaCore_718

//KaratsubaCore_366 replaced by KaratsubaCore_717

//BADD_999 replaced by BADD_1412

//BADD_998 replaced by BADD_1411

//BADD_997 replaced by BADD_1410

//KaratsubaCore_371 replaced by KaratsubaCore_717

//KaratsubaCore_370 replaced by KaratsubaCore_718

//KaratsubaCore_369 replaced by KaratsubaCore_717

//BADD_1003 replaced by BADD_1406

//BADD_1002 replaced by BADD_1408

//BADD_1001 replaced by BADD_1407

//BADD_1000 replaced by BADD_1406

//KaratsubaCore_374 replaced by KaratsubaCore_718

//KaratsubaCore_373 replaced by KaratsubaCore_715

//KaratsubaCore_372 replaced by KaratsubaCore_718

//BADD_1006 replaced by BADD_1412

//BADD_1005 replaced by BADD_1411

//BADD_1004 replaced by BADD_1410

//KaratsubaCore_377 replaced by KaratsubaCore_717

//KaratsubaCore_376 replaced by KaratsubaCore_718

//KaratsubaCore_375 replaced by KaratsubaCore_717

//BADD_1010 replaced by BADD_1406

//BADD_1009 replaced by BADD_1408

//BADD_1008 replaced by BADD_1407

//BADD_1007 replaced by BADD_1406

//KaratsubaCore_380 replaced by KaratsubaCore_718

//KaratsubaCore_379 replaced by KaratsubaCore_715

//KaratsubaCore_378 replaced by KaratsubaCore_718

//BADD_1014 replaced by BADD_1395

//BADD_1013 replaced by BADD_1397

//BADD_1012 replaced by BADD_1396

//BADD_1011 replaced by BADD_1395

//KaratsubaCore_383 replaced by KaratsubaCore_715

//KaratsubaCore_382 replaced by KaratsubaCore_706

//KaratsubaCore_381 replaced by KaratsubaCore_715

//BADD_1018 replaced by BADD_1406

//BADD_1017 replaced by BADD_1408

//BADD_1016 replaced by BADD_1407

//BADD_1015 replaced by BADD_1406

//KaratsubaCore_386 replaced by KaratsubaCore_718

//KaratsubaCore_385 replaced by KaratsubaCore_715

//KaratsubaCore_384 replaced by KaratsubaCore_718

//BADD_1021 replaced by BADD_1412

//BADD_1020 replaced by BADD_1411

//BADD_1019 replaced by BADD_1410

//KaratsubaCore_389 replaced by KaratsubaCore_717

//KaratsubaCore_388 replaced by KaratsubaCore_718

//KaratsubaCore_387 replaced by KaratsubaCore_717

//BADD_1025 replaced by BADD_1406

//BADD_1024 replaced by BADD_1408

//BADD_1023 replaced by BADD_1407

//BADD_1022 replaced by BADD_1406

//KaratsubaCore_392 replaced by KaratsubaCore_718

//KaratsubaCore_391 replaced by KaratsubaCore_715

//KaratsubaCore_390 replaced by KaratsubaCore_718

//BADD_1028 replaced by BADD_1412

//BADD_1027 replaced by BADD_1411

//BADD_1026 replaced by BADD_1410

//KaratsubaCore_395 replaced by KaratsubaCore_717

//KaratsubaCore_394 replaced by KaratsubaCore_718

//KaratsubaCore_393 replaced by KaratsubaCore_717

//BADD_1031 replaced by BADD_1412

//BADD_1030 replaced by BADD_1411

//BADD_1029 replaced by BADD_1410

//KaratsubaCore_398 replaced by KaratsubaCore_717

//KaratsubaCore_397 replaced by KaratsubaCore_718

//KaratsubaCore_396 replaced by KaratsubaCore_717

//BADD_1035 replaced by BADD_1406

//BADD_1034 replaced by BADD_1408

//BADD_1033 replaced by BADD_1407

//BADD_1032 replaced by BADD_1406

//KaratsubaCore_401 replaced by KaratsubaCore_718

//KaratsubaCore_400 replaced by KaratsubaCore_715

//KaratsubaCore_399 replaced by KaratsubaCore_718

//BADD_1038 replaced by BADD_1412

//BADD_1037 replaced by BADD_1411

//BADD_1036 replaced by BADD_1410

//KaratsubaCore_404 replaced by KaratsubaCore_717

//KaratsubaCore_403 replaced by KaratsubaCore_718

//KaratsubaCore_402 replaced by KaratsubaCore_717

//BADD_1042 replaced by BADD_1406

//BADD_1041 replaced by BADD_1408

//BADD_1040 replaced by BADD_1407

//BADD_1039 replaced by BADD_1406

//KaratsubaCore_407 replaced by KaratsubaCore_718

//KaratsubaCore_406 replaced by KaratsubaCore_715

//KaratsubaCore_405 replaced by KaratsubaCore_718

//BADD_1046 replaced by BADD_1395

//BADD_1045 replaced by BADD_1397

//BADD_1044 replaced by BADD_1396

//BADD_1043 replaced by BADD_1395

//KaratsubaCore_410 replaced by KaratsubaCore_715

//KaratsubaCore_409 replaced by KaratsubaCore_706

//KaratsubaCore_408 replaced by KaratsubaCore_715

//BADD_1050 replaced by BADD_1406

//BADD_1049 replaced by BADD_1408

//BADD_1048 replaced by BADD_1407

//BADD_1047 replaced by BADD_1406

//KaratsubaCore_413 replaced by KaratsubaCore_718

//KaratsubaCore_412 replaced by KaratsubaCore_715

//KaratsubaCore_411 replaced by KaratsubaCore_718

//BADD_1053 replaced by BADD_1412

//BADD_1052 replaced by BADD_1411

//BADD_1051 replaced by BADD_1410

//KaratsubaCore_416 replaced by KaratsubaCore_717

//KaratsubaCore_415 replaced by KaratsubaCore_718

//KaratsubaCore_414 replaced by KaratsubaCore_717

//BADD_1057 replaced by BADD_1406

//BADD_1056 replaced by BADD_1408

//BADD_1055 replaced by BADD_1407

//BADD_1054 replaced by BADD_1406

//KaratsubaCore_419 replaced by KaratsubaCore_718

//KaratsubaCore_418 replaced by KaratsubaCore_715

//KaratsubaCore_417 replaced by KaratsubaCore_718

//BADD_1060 replaced by BADD_1412

//BADD_1059 replaced by BADD_1411

//BADD_1058 replaced by BADD_1410

//KaratsubaCore_422 replaced by KaratsubaCore_717

//KaratsubaCore_421 replaced by KaratsubaCore_718

//KaratsubaCore_420 replaced by KaratsubaCore_717

//BADD_1063 replaced by BADD_1412

//BADD_1062 replaced by BADD_1411

//BADD_1061 replaced by BADD_1410

//KaratsubaCore_425 replaced by KaratsubaCore_717

//KaratsubaCore_424 replaced by KaratsubaCore_718

//KaratsubaCore_423 replaced by KaratsubaCore_717

//BADD_1067 replaced by BADD_1406

//BADD_1066 replaced by BADD_1408

//BADD_1065 replaced by BADD_1407

//BADD_1064 replaced by BADD_1406

//KaratsubaCore_428 replaced by KaratsubaCore_718

//KaratsubaCore_427 replaced by KaratsubaCore_715

//KaratsubaCore_426 replaced by KaratsubaCore_718

//BADD_1070 replaced by BADD_1412

//BADD_1069 replaced by BADD_1411

//BADD_1068 replaced by BADD_1410

//KaratsubaCore_431 replaced by KaratsubaCore_717

//KaratsubaCore_430 replaced by KaratsubaCore_718

//KaratsubaCore_429 replaced by KaratsubaCore_717

//BADD_1074 replaced by BADD_1406

//BADD_1073 replaced by BADD_1408

//BADD_1072 replaced by BADD_1407

//BADD_1071 replaced by BADD_1406

//KaratsubaCore_434 replaced by KaratsubaCore_718

//KaratsubaCore_433 replaced by KaratsubaCore_715

//KaratsubaCore_432 replaced by KaratsubaCore_718

//BADD_1078 replaced by BADD_1395

//BADD_1077 replaced by BADD_1397

//BADD_1076 replaced by BADD_1396

//BADD_1075 replaced by BADD_1395

//KaratsubaCore_437 replaced by KaratsubaCore_715

//KaratsubaCore_436 replaced by KaratsubaCore_706

//KaratsubaCore_435 replaced by KaratsubaCore_715

//BADD_1082 replaced by BADD_1406

//BADD_1081 replaced by BADD_1408

//BADD_1080 replaced by BADD_1407

//BADD_1079 replaced by BADD_1406

//KaratsubaCore_440 replaced by KaratsubaCore_718

//KaratsubaCore_439 replaced by KaratsubaCore_715

//KaratsubaCore_438 replaced by KaratsubaCore_718

//BADD_1085 replaced by BADD_1412

//BADD_1084 replaced by BADD_1411

//BADD_1083 replaced by BADD_1410

//KaratsubaCore_443 replaced by KaratsubaCore_717

//KaratsubaCore_442 replaced by KaratsubaCore_718

//KaratsubaCore_441 replaced by KaratsubaCore_717

//BADD_1089 replaced by BADD_1406

//BADD_1088 replaced by BADD_1408

//BADD_1087 replaced by BADD_1407

//BADD_1086 replaced by BADD_1406

//KaratsubaCore_446 replaced by KaratsubaCore_718

//KaratsubaCore_445 replaced by KaratsubaCore_715

//KaratsubaCore_444 replaced by KaratsubaCore_718

//BADD_1092 replaced by BADD_1412

//BADD_1091 replaced by BADD_1411

//BADD_1090 replaced by BADD_1410

//KaratsubaCore_449 replaced by KaratsubaCore_717

//KaratsubaCore_448 replaced by KaratsubaCore_718

//KaratsubaCore_447 replaced by KaratsubaCore_717

//BADD_1095 replaced by BADD_1412

//BADD_1094 replaced by BADD_1411

//BADD_1093 replaced by BADD_1410

//KaratsubaCore_452 replaced by KaratsubaCore_717

//KaratsubaCore_451 replaced by KaratsubaCore_718

//KaratsubaCore_450 replaced by KaratsubaCore_717

//BADD_1099 replaced by BADD_1406

//BADD_1098 replaced by BADD_1408

//BADD_1097 replaced by BADD_1407

//BADD_1096 replaced by BADD_1406

//KaratsubaCore_455 replaced by KaratsubaCore_718

//KaratsubaCore_454 replaced by KaratsubaCore_715

//KaratsubaCore_453 replaced by KaratsubaCore_718

//BADD_1102 replaced by BADD_1412

//BADD_1101 replaced by BADD_1411

//BADD_1100 replaced by BADD_1410

//KaratsubaCore_458 replaced by KaratsubaCore_717

//KaratsubaCore_457 replaced by KaratsubaCore_718

//KaratsubaCore_456 replaced by KaratsubaCore_717

//BADD_1106 replaced by BADD_1406

//BADD_1105 replaced by BADD_1408

//BADD_1104 replaced by BADD_1407

//BADD_1103 replaced by BADD_1406

//KaratsubaCore_461 replaced by KaratsubaCore_718

//KaratsubaCore_460 replaced by KaratsubaCore_715

//KaratsubaCore_459 replaced by KaratsubaCore_718

//BADD_1110 replaced by BADD_1395

//BADD_1109 replaced by BADD_1397

//BADD_1108 replaced by BADD_1396

//BADD_1107 replaced by BADD_1395

//KaratsubaCore_464 replaced by KaratsubaCore_715

//KaratsubaCore_463 replaced by KaratsubaCore_706

//KaratsubaCore_462 replaced by KaratsubaCore_715

//BADD_1114 replaced by BADD_1406

//BADD_1113 replaced by BADD_1408

//BADD_1112 replaced by BADD_1407

//BADD_1111 replaced by BADD_1406

//KaratsubaCore_467 replaced by KaratsubaCore_718

//KaratsubaCore_466 replaced by KaratsubaCore_715

//KaratsubaCore_465 replaced by KaratsubaCore_718

//BADD_1117 replaced by BADD_1412

//BADD_1116 replaced by BADD_1411

//BADD_1115 replaced by BADD_1410

//KaratsubaCore_470 replaced by KaratsubaCore_717

//KaratsubaCore_469 replaced by KaratsubaCore_718

//KaratsubaCore_468 replaced by KaratsubaCore_717

//BADD_1121 replaced by BADD_1406

//BADD_1120 replaced by BADD_1408

//BADD_1119 replaced by BADD_1407

//BADD_1118 replaced by BADD_1406

//KaratsubaCore_473 replaced by KaratsubaCore_718

//KaratsubaCore_472 replaced by KaratsubaCore_715

//KaratsubaCore_471 replaced by KaratsubaCore_718

//BADD_1124 replaced by BADD_1412

//BADD_1123 replaced by BADD_1411

//BADD_1122 replaced by BADD_1410

//KaratsubaCore_476 replaced by KaratsubaCore_717

//KaratsubaCore_475 replaced by KaratsubaCore_718

//KaratsubaCore_474 replaced by KaratsubaCore_717

//BADD_1127 replaced by BADD_1412

//BADD_1126 replaced by BADD_1411

//BADD_1125 replaced by BADD_1410

//KaratsubaCore_479 replaced by KaratsubaCore_717

//KaratsubaCore_478 replaced by KaratsubaCore_718

//KaratsubaCore_477 replaced by KaratsubaCore_717

//BADD_1131 replaced by BADD_1406

//BADD_1130 replaced by BADD_1408

//BADD_1129 replaced by BADD_1407

//BADD_1128 replaced by BADD_1406

//KaratsubaCore_482 replaced by KaratsubaCore_718

//KaratsubaCore_481 replaced by KaratsubaCore_715

//KaratsubaCore_480 replaced by KaratsubaCore_718

//BADD_1134 replaced by BADD_1412

//BADD_1133 replaced by BADD_1411

//BADD_1132 replaced by BADD_1410

//KaratsubaCore_485 replaced by KaratsubaCore_717

//KaratsubaCore_484 replaced by KaratsubaCore_718

//KaratsubaCore_483 replaced by KaratsubaCore_717

//BADD_1138 replaced by BADD_1406

//BADD_1137 replaced by BADD_1408

//BADD_1136 replaced by BADD_1407

//BADD_1135 replaced by BADD_1406

//KaratsubaCore_488 replaced by KaratsubaCore_718

//KaratsubaCore_487 replaced by KaratsubaCore_715

//KaratsubaCore_486 replaced by KaratsubaCore_718

//BADD_1142 replaced by BADD_1395

//BADD_1141 replaced by BADD_1397

//BADD_1140 replaced by BADD_1396

//BADD_1139 replaced by BADD_1395

//KaratsubaCore_491 replaced by KaratsubaCore_715

//KaratsubaCore_490 replaced by KaratsubaCore_706

//KaratsubaCore_489 replaced by KaratsubaCore_715

//BADD_1146 replaced by BADD_1406

//BADD_1145 replaced by BADD_1408

//BADD_1144 replaced by BADD_1407

//BADD_1143 replaced by BADD_1406

//KaratsubaCore_494 replaced by KaratsubaCore_718

//KaratsubaCore_493 replaced by KaratsubaCore_715

//KaratsubaCore_492 replaced by KaratsubaCore_718

//BADD_1149 replaced by BADD_1412

//BADD_1148 replaced by BADD_1411

//BADD_1147 replaced by BADD_1410

//KaratsubaCore_497 replaced by KaratsubaCore_717

//KaratsubaCore_496 replaced by KaratsubaCore_718

//KaratsubaCore_495 replaced by KaratsubaCore_717

//BADD_1153 replaced by BADD_1406

//BADD_1152 replaced by BADD_1408

//BADD_1151 replaced by BADD_1407

//BADD_1150 replaced by BADD_1406

//KaratsubaCore_500 replaced by KaratsubaCore_718

//KaratsubaCore_499 replaced by KaratsubaCore_715

//KaratsubaCore_498 replaced by KaratsubaCore_718

//BADD_1156 replaced by BADD_1412

//BADD_1155 replaced by BADD_1411

//BADD_1154 replaced by BADD_1410

//KaratsubaCore_503 replaced by KaratsubaCore_717

//KaratsubaCore_502 replaced by KaratsubaCore_718

//KaratsubaCore_501 replaced by KaratsubaCore_717

//BADD_1159 replaced by BADD_1412

//BADD_1158 replaced by BADD_1411

//BADD_1157 replaced by BADD_1410

//KaratsubaCore_506 replaced by KaratsubaCore_717

//KaratsubaCore_505 replaced by KaratsubaCore_718

//KaratsubaCore_504 replaced by KaratsubaCore_717

//BADD_1163 replaced by BADD_1406

//BADD_1162 replaced by BADD_1408

//BADD_1161 replaced by BADD_1407

//BADD_1160 replaced by BADD_1406

//KaratsubaCore_509 replaced by KaratsubaCore_718

//KaratsubaCore_508 replaced by KaratsubaCore_715

//KaratsubaCore_507 replaced by KaratsubaCore_718

//BADD_1166 replaced by BADD_1412

//BADD_1165 replaced by BADD_1411

//BADD_1164 replaced by BADD_1410

//KaratsubaCore_512 replaced by KaratsubaCore_717

//KaratsubaCore_511 replaced by KaratsubaCore_718

//KaratsubaCore_510 replaced by KaratsubaCore_717

//BADD_1170 replaced by BADD_1406

//BADD_1169 replaced by BADD_1408

//BADD_1168 replaced by BADD_1407

//BADD_1167 replaced by BADD_1406

//KaratsubaCore_515 replaced by KaratsubaCore_718

//KaratsubaCore_514 replaced by KaratsubaCore_715

//KaratsubaCore_513 replaced by KaratsubaCore_718

//BADD_1174 replaced by BADD_1395

//BADD_1173 replaced by BADD_1397

//BADD_1172 replaced by BADD_1396

//BADD_1171 replaced by BADD_1395

//KaratsubaCore_518 replaced by KaratsubaCore_715

//KaratsubaCore_517 replaced by KaratsubaCore_706

//KaratsubaCore_516 replaced by KaratsubaCore_715

//BADD_1178 replaced by BADD_1406

//BADD_1177 replaced by BADD_1408

//BADD_1176 replaced by BADD_1407

//BADD_1175 replaced by BADD_1406

//KaratsubaCore_521 replaced by KaratsubaCore_718

//KaratsubaCore_520 replaced by KaratsubaCore_715

//KaratsubaCore_519 replaced by KaratsubaCore_718

//BADD_1181 replaced by BADD_1412

//BADD_1180 replaced by BADD_1411

//BADD_1179 replaced by BADD_1410

//KaratsubaCore_524 replaced by KaratsubaCore_717

//KaratsubaCore_523 replaced by KaratsubaCore_718

//KaratsubaCore_522 replaced by KaratsubaCore_717

//BADD_1185 replaced by BADD_1406

//BADD_1184 replaced by BADD_1408

//BADD_1183 replaced by BADD_1407

//BADD_1182 replaced by BADD_1406

//KaratsubaCore_527 replaced by KaratsubaCore_718

//KaratsubaCore_526 replaced by KaratsubaCore_715

//KaratsubaCore_525 replaced by KaratsubaCore_718

//BADD_1188 replaced by BADD_1412

//BADD_1187 replaced by BADD_1411

//BADD_1186 replaced by BADD_1410

//KaratsubaCore_530 replaced by KaratsubaCore_717

//KaratsubaCore_529 replaced by KaratsubaCore_718

//KaratsubaCore_528 replaced by KaratsubaCore_717

//BADD_1191 replaced by BADD_1412

//BADD_1190 replaced by BADD_1411

//BADD_1189 replaced by BADD_1410

//KaratsubaCore_533 replaced by KaratsubaCore_717

//KaratsubaCore_532 replaced by KaratsubaCore_718

//KaratsubaCore_531 replaced by KaratsubaCore_717

//BADD_1195 replaced by BADD_1406

//BADD_1194 replaced by BADD_1408

//BADD_1193 replaced by BADD_1407

//BADD_1192 replaced by BADD_1406

//KaratsubaCore_536 replaced by KaratsubaCore_718

//KaratsubaCore_535 replaced by KaratsubaCore_715

//KaratsubaCore_534 replaced by KaratsubaCore_718

//BADD_1198 replaced by BADD_1412

//BADD_1197 replaced by BADD_1411

//BADD_1196 replaced by BADD_1410

//KaratsubaCore_539 replaced by KaratsubaCore_717

//KaratsubaCore_538 replaced by KaratsubaCore_718

//KaratsubaCore_537 replaced by KaratsubaCore_717

//BADD_1202 replaced by BADD_1406

//BADD_1201 replaced by BADD_1408

//BADD_1200 replaced by BADD_1407

//BADD_1199 replaced by BADD_1406

//KaratsubaCore_542 replaced by KaratsubaCore_718

//KaratsubaCore_541 replaced by KaratsubaCore_715

//KaratsubaCore_540 replaced by KaratsubaCore_718

//BADD_1206 replaced by BADD_1395

//BADD_1205 replaced by BADD_1397

//BADD_1204 replaced by BADD_1396

//BADD_1203 replaced by BADD_1395

//KaratsubaCore_545 replaced by KaratsubaCore_715

//KaratsubaCore_544 replaced by KaratsubaCore_706

//KaratsubaCore_543 replaced by KaratsubaCore_715

//BADD_1210 replaced by BADD_1406

//BADD_1209 replaced by BADD_1408

//BADD_1208 replaced by BADD_1407

//BADD_1207 replaced by BADD_1406

//KaratsubaCore_548 replaced by KaratsubaCore_718

//KaratsubaCore_547 replaced by KaratsubaCore_715

//KaratsubaCore_546 replaced by KaratsubaCore_718

//BADD_1213 replaced by BADD_1412

//BADD_1212 replaced by BADD_1411

//BADD_1211 replaced by BADD_1410

//KaratsubaCore_551 replaced by KaratsubaCore_717

//KaratsubaCore_550 replaced by KaratsubaCore_718

//KaratsubaCore_549 replaced by KaratsubaCore_717

//BADD_1217 replaced by BADD_1406

//BADD_1216 replaced by BADD_1408

//BADD_1215 replaced by BADD_1407

//BADD_1214 replaced by BADD_1406

//KaratsubaCore_554 replaced by KaratsubaCore_718

//KaratsubaCore_553 replaced by KaratsubaCore_715

//KaratsubaCore_552 replaced by KaratsubaCore_718

//BADD_1220 replaced by BADD_1412

//BADD_1219 replaced by BADD_1411

//BADD_1218 replaced by BADD_1410

//KaratsubaCore_557 replaced by KaratsubaCore_717

//KaratsubaCore_556 replaced by KaratsubaCore_718

//KaratsubaCore_555 replaced by KaratsubaCore_717

//BADD_1223 replaced by BADD_1412

//BADD_1222 replaced by BADD_1411

//BADD_1221 replaced by BADD_1410

//KaratsubaCore_560 replaced by KaratsubaCore_717

//KaratsubaCore_559 replaced by KaratsubaCore_718

//KaratsubaCore_558 replaced by KaratsubaCore_717

//BADD_1227 replaced by BADD_1406

//BADD_1226 replaced by BADD_1408

//BADD_1225 replaced by BADD_1407

//BADD_1224 replaced by BADD_1406

//KaratsubaCore_563 replaced by KaratsubaCore_718

//KaratsubaCore_562 replaced by KaratsubaCore_715

//KaratsubaCore_561 replaced by KaratsubaCore_718

//BADD_1230 replaced by BADD_1412

//BADD_1229 replaced by BADD_1411

//BADD_1228 replaced by BADD_1410

//KaratsubaCore_566 replaced by KaratsubaCore_717

//KaratsubaCore_565 replaced by KaratsubaCore_718

//KaratsubaCore_564 replaced by KaratsubaCore_717

//BADD_1234 replaced by BADD_1406

//BADD_1233 replaced by BADD_1408

//BADD_1232 replaced by BADD_1407

//BADD_1231 replaced by BADD_1406

//KaratsubaCore_569 replaced by KaratsubaCore_718

//KaratsubaCore_568 replaced by KaratsubaCore_715

//KaratsubaCore_567 replaced by KaratsubaCore_718

//BADD_1238 replaced by BADD_1395

//BADD_1237 replaced by BADD_1397

//BADD_1236 replaced by BADD_1396

//BADD_1235 replaced by BADD_1395

//KaratsubaCore_572 replaced by KaratsubaCore_715

//KaratsubaCore_571 replaced by KaratsubaCore_706

//KaratsubaCore_570 replaced by KaratsubaCore_715

//BADD_1242 replaced by BADD_1406

//BADD_1241 replaced by BADD_1408

//BADD_1240 replaced by BADD_1407

//BADD_1239 replaced by BADD_1406

//KaratsubaCore_575 replaced by KaratsubaCore_718

//KaratsubaCore_574 replaced by KaratsubaCore_715

//KaratsubaCore_573 replaced by KaratsubaCore_718

//BADD_1245 replaced by BADD_1412

//BADD_1244 replaced by BADD_1411

//BADD_1243 replaced by BADD_1410

//KaratsubaCore_578 replaced by KaratsubaCore_717

//KaratsubaCore_577 replaced by KaratsubaCore_718

//KaratsubaCore_576 replaced by KaratsubaCore_717

//BADD_1249 replaced by BADD_1406

//BADD_1248 replaced by BADD_1408

//BADD_1247 replaced by BADD_1407

//BADD_1246 replaced by BADD_1406

//KaratsubaCore_581 replaced by KaratsubaCore_718

//KaratsubaCore_580 replaced by KaratsubaCore_715

//KaratsubaCore_579 replaced by KaratsubaCore_718

//BADD_1252 replaced by BADD_1412

//BADD_1251 replaced by BADD_1411

//BADD_1250 replaced by BADD_1410

//KaratsubaCore_584 replaced by KaratsubaCore_717

//KaratsubaCore_583 replaced by KaratsubaCore_718

//KaratsubaCore_582 replaced by KaratsubaCore_717

//BADD_1255 replaced by BADD_1412

//BADD_1254 replaced by BADD_1411

//BADD_1253 replaced by BADD_1410

//KaratsubaCore_587 replaced by KaratsubaCore_717

//KaratsubaCore_586 replaced by KaratsubaCore_718

//KaratsubaCore_585 replaced by KaratsubaCore_717

//BADD_1259 replaced by BADD_1406

//BADD_1258 replaced by BADD_1408

//BADD_1257 replaced by BADD_1407

//BADD_1256 replaced by BADD_1406

//KaratsubaCore_590 replaced by KaratsubaCore_718

//KaratsubaCore_589 replaced by KaratsubaCore_715

//KaratsubaCore_588 replaced by KaratsubaCore_718

//BADD_1262 replaced by BADD_1412

//BADD_1261 replaced by BADD_1411

//BADD_1260 replaced by BADD_1410

//KaratsubaCore_593 replaced by KaratsubaCore_717

//KaratsubaCore_592 replaced by KaratsubaCore_718

//KaratsubaCore_591 replaced by KaratsubaCore_717

//BADD_1266 replaced by BADD_1406

//BADD_1265 replaced by BADD_1408

//BADD_1264 replaced by BADD_1407

//BADD_1263 replaced by BADD_1406

//KaratsubaCore_596 replaced by KaratsubaCore_718

//KaratsubaCore_595 replaced by KaratsubaCore_715

//KaratsubaCore_594 replaced by KaratsubaCore_718

//BADD_1270 replaced by BADD_1395

//BADD_1269 replaced by BADD_1397

//BADD_1268 replaced by BADD_1396

//BADD_1267 replaced by BADD_1395

//KaratsubaCore_599 replaced by KaratsubaCore_715

//KaratsubaCore_598 replaced by KaratsubaCore_706

//KaratsubaCore_597 replaced by KaratsubaCore_715

//BADD_1274 replaced by BADD_1406

//BADD_1273 replaced by BADD_1408

//BADD_1272 replaced by BADD_1407

//BADD_1271 replaced by BADD_1406

//KaratsubaCore_602 replaced by KaratsubaCore_718

//KaratsubaCore_601 replaced by KaratsubaCore_715

//KaratsubaCore_600 replaced by KaratsubaCore_718

//BADD_1277 replaced by BADD_1412

//BADD_1276 replaced by BADD_1411

//BADD_1275 replaced by BADD_1410

//KaratsubaCore_605 replaced by KaratsubaCore_717

//KaratsubaCore_604 replaced by KaratsubaCore_718

//KaratsubaCore_603 replaced by KaratsubaCore_717

//BADD_1281 replaced by BADD_1406

//BADD_1280 replaced by BADD_1408

//BADD_1279 replaced by BADD_1407

//BADD_1278 replaced by BADD_1406

//KaratsubaCore_608 replaced by KaratsubaCore_718

//KaratsubaCore_607 replaced by KaratsubaCore_715

//KaratsubaCore_606 replaced by KaratsubaCore_718

//BADD_1284 replaced by BADD_1412

//BADD_1283 replaced by BADD_1411

//BADD_1282 replaced by BADD_1410

//KaratsubaCore_611 replaced by KaratsubaCore_717

//KaratsubaCore_610 replaced by KaratsubaCore_718

//KaratsubaCore_609 replaced by KaratsubaCore_717

//BADD_1287 replaced by BADD_1412

//BADD_1286 replaced by BADD_1411

//BADD_1285 replaced by BADD_1410

//KaratsubaCore_614 replaced by KaratsubaCore_717

//KaratsubaCore_613 replaced by KaratsubaCore_718

//KaratsubaCore_612 replaced by KaratsubaCore_717

//BADD_1291 replaced by BADD_1406

//BADD_1290 replaced by BADD_1408

//BADD_1289 replaced by BADD_1407

//BADD_1288 replaced by BADD_1406

//KaratsubaCore_617 replaced by KaratsubaCore_718

//KaratsubaCore_616 replaced by KaratsubaCore_715

//KaratsubaCore_615 replaced by KaratsubaCore_718

//BADD_1294 replaced by BADD_1412

//BADD_1293 replaced by BADD_1411

//BADD_1292 replaced by BADD_1410

//KaratsubaCore_620 replaced by KaratsubaCore_717

//KaratsubaCore_619 replaced by KaratsubaCore_718

//KaratsubaCore_618 replaced by KaratsubaCore_717

//BADD_1298 replaced by BADD_1406

//BADD_1297 replaced by BADD_1408

//BADD_1296 replaced by BADD_1407

//BADD_1295 replaced by BADD_1406

//KaratsubaCore_623 replaced by KaratsubaCore_718

//KaratsubaCore_622 replaced by KaratsubaCore_715

//KaratsubaCore_621 replaced by KaratsubaCore_718

//BADD_1302 replaced by BADD_1395

//BADD_1301 replaced by BADD_1397

//BADD_1300 replaced by BADD_1396

//BADD_1299 replaced by BADD_1395

//KaratsubaCore_626 replaced by KaratsubaCore_715

//KaratsubaCore_625 replaced by KaratsubaCore_706

//KaratsubaCore_624 replaced by KaratsubaCore_715

//BADD_1306 replaced by BADD_1406

//BADD_1305 replaced by BADD_1408

//BADD_1304 replaced by BADD_1407

//BADD_1303 replaced by BADD_1406

//KaratsubaCore_629 replaced by KaratsubaCore_718

//KaratsubaCore_628 replaced by KaratsubaCore_715

//KaratsubaCore_627 replaced by KaratsubaCore_718

//BADD_1309 replaced by BADD_1412

//BADD_1308 replaced by BADD_1411

//BADD_1307 replaced by BADD_1410

//KaratsubaCore_632 replaced by KaratsubaCore_717

//KaratsubaCore_631 replaced by KaratsubaCore_718

//KaratsubaCore_630 replaced by KaratsubaCore_717

//BADD_1313 replaced by BADD_1406

//BADD_1312 replaced by BADD_1408

//BADD_1311 replaced by BADD_1407

//BADD_1310 replaced by BADD_1406

//KaratsubaCore_635 replaced by KaratsubaCore_718

//KaratsubaCore_634 replaced by KaratsubaCore_715

//KaratsubaCore_633 replaced by KaratsubaCore_718

//BADD_1316 replaced by BADD_1412

//BADD_1315 replaced by BADD_1411

//BADD_1314 replaced by BADD_1410

//KaratsubaCore_638 replaced by KaratsubaCore_717

//KaratsubaCore_637 replaced by KaratsubaCore_718

//KaratsubaCore_636 replaced by KaratsubaCore_717

//BADD_1319 replaced by BADD_1412

//BADD_1318 replaced by BADD_1411

//BADD_1317 replaced by BADD_1410

//KaratsubaCore_641 replaced by KaratsubaCore_717

//KaratsubaCore_640 replaced by KaratsubaCore_718

//KaratsubaCore_639 replaced by KaratsubaCore_717

//BADD_1323 replaced by BADD_1406

//BADD_1322 replaced by BADD_1408

//BADD_1321 replaced by BADD_1407

//BADD_1320 replaced by BADD_1406

//KaratsubaCore_644 replaced by KaratsubaCore_718

//KaratsubaCore_643 replaced by KaratsubaCore_715

//KaratsubaCore_642 replaced by KaratsubaCore_718

//BADD_1326 replaced by BADD_1412

//BADD_1325 replaced by BADD_1411

//BADD_1324 replaced by BADD_1410

//KaratsubaCore_647 replaced by KaratsubaCore_717

//KaratsubaCore_646 replaced by KaratsubaCore_718

//KaratsubaCore_645 replaced by KaratsubaCore_717

//BADD_1330 replaced by BADD_1406

//BADD_1329 replaced by BADD_1408

//BADD_1328 replaced by BADD_1407

//BADD_1327 replaced by BADD_1406

//KaratsubaCore_650 replaced by KaratsubaCore_718

//KaratsubaCore_649 replaced by KaratsubaCore_715

//KaratsubaCore_648 replaced by KaratsubaCore_718

//BADD_1334 replaced by BADD_1395

//BADD_1333 replaced by BADD_1397

//BADD_1332 replaced by BADD_1396

//BADD_1331 replaced by BADD_1395

//KaratsubaCore_653 replaced by KaratsubaCore_715

//KaratsubaCore_652 replaced by KaratsubaCore_706

//KaratsubaCore_651 replaced by KaratsubaCore_715

//BADD_1338 replaced by BADD_1406

//BADD_1337 replaced by BADD_1408

//BADD_1336 replaced by BADD_1407

//BADD_1335 replaced by BADD_1406

//KaratsubaCore_656 replaced by KaratsubaCore_718

//KaratsubaCore_655 replaced by KaratsubaCore_715

//KaratsubaCore_654 replaced by KaratsubaCore_718

//BADD_1341 replaced by BADD_1412

//BADD_1340 replaced by BADD_1411

//BADD_1339 replaced by BADD_1410

//KaratsubaCore_659 replaced by KaratsubaCore_717

//KaratsubaCore_658 replaced by KaratsubaCore_718

//KaratsubaCore_657 replaced by KaratsubaCore_717

//BADD_1345 replaced by BADD_1406

//BADD_1344 replaced by BADD_1408

//BADD_1343 replaced by BADD_1407

//BADD_1342 replaced by BADD_1406

//KaratsubaCore_662 replaced by KaratsubaCore_718

//KaratsubaCore_661 replaced by KaratsubaCore_715

//KaratsubaCore_660 replaced by KaratsubaCore_718

//BADD_1348 replaced by BADD_1412

//BADD_1347 replaced by BADD_1411

//BADD_1346 replaced by BADD_1410

//KaratsubaCore_665 replaced by KaratsubaCore_717

//KaratsubaCore_664 replaced by KaratsubaCore_718

//KaratsubaCore_663 replaced by KaratsubaCore_717

//BADD_1351 replaced by BADD_1412

//BADD_1350 replaced by BADD_1411

//BADD_1349 replaced by BADD_1410

//KaratsubaCore_668 replaced by KaratsubaCore_717

//KaratsubaCore_667 replaced by KaratsubaCore_718

//KaratsubaCore_666 replaced by KaratsubaCore_717

//BADD_1355 replaced by BADD_1406

//BADD_1354 replaced by BADD_1408

//BADD_1353 replaced by BADD_1407

//BADD_1352 replaced by BADD_1406

//KaratsubaCore_671 replaced by KaratsubaCore_718

//KaratsubaCore_670 replaced by KaratsubaCore_715

//KaratsubaCore_669 replaced by KaratsubaCore_718

//BADD_1358 replaced by BADD_1412

//BADD_1357 replaced by BADD_1411

//BADD_1356 replaced by BADD_1410

//KaratsubaCore_674 replaced by KaratsubaCore_717

//KaratsubaCore_673 replaced by KaratsubaCore_718

//KaratsubaCore_672 replaced by KaratsubaCore_717

//BADD_1362 replaced by BADD_1406

//BADD_1361 replaced by BADD_1408

//BADD_1360 replaced by BADD_1407

//BADD_1359 replaced by BADD_1406

//KaratsubaCore_677 replaced by KaratsubaCore_718

//KaratsubaCore_676 replaced by KaratsubaCore_715

//KaratsubaCore_675 replaced by KaratsubaCore_718

//BADD_1366 replaced by BADD_1395

//BADD_1365 replaced by BADD_1397

//BADD_1364 replaced by BADD_1396

//BADD_1363 replaced by BADD_1395

//KaratsubaCore_680 replaced by KaratsubaCore_715

//KaratsubaCore_679 replaced by KaratsubaCore_706

//KaratsubaCore_678 replaced by KaratsubaCore_715

//BADD_1370 replaced by BADD_1406

//BADD_1369 replaced by BADD_1408

//BADD_1368 replaced by BADD_1407

//BADD_1367 replaced by BADD_1406

//KaratsubaCore_683 replaced by KaratsubaCore_718

//KaratsubaCore_682 replaced by KaratsubaCore_715

//KaratsubaCore_681 replaced by KaratsubaCore_718

//BADD_1373 replaced by BADD_1412

//BADD_1372 replaced by BADD_1411

//BADD_1371 replaced by BADD_1410

//KaratsubaCore_686 replaced by KaratsubaCore_717

//KaratsubaCore_685 replaced by KaratsubaCore_718

//KaratsubaCore_684 replaced by KaratsubaCore_717

//BADD_1377 replaced by BADD_1406

//BADD_1376 replaced by BADD_1408

//BADD_1375 replaced by BADD_1407

//BADD_1374 replaced by BADD_1406

//KaratsubaCore_689 replaced by KaratsubaCore_718

//KaratsubaCore_688 replaced by KaratsubaCore_715

//KaratsubaCore_687 replaced by KaratsubaCore_718

//BADD_1380 replaced by BADD_1412

//BADD_1379 replaced by BADD_1411

//BADD_1378 replaced by BADD_1410

//KaratsubaCore_692 replaced by KaratsubaCore_717

//KaratsubaCore_691 replaced by KaratsubaCore_718

//KaratsubaCore_690 replaced by KaratsubaCore_717

//BADD_1383 replaced by BADD_1412

//BADD_1382 replaced by BADD_1411

//BADD_1381 replaced by BADD_1410

//KaratsubaCore_695 replaced by KaratsubaCore_717

//KaratsubaCore_694 replaced by KaratsubaCore_718

//KaratsubaCore_693 replaced by KaratsubaCore_717

//BADD_1387 replaced by BADD_1406

//BADD_1386 replaced by BADD_1408

//BADD_1385 replaced by BADD_1407

//BADD_1384 replaced by BADD_1406

//KaratsubaCore_698 replaced by KaratsubaCore_718

//KaratsubaCore_697 replaced by KaratsubaCore_715

//KaratsubaCore_696 replaced by KaratsubaCore_718

//BADD_1390 replaced by BADD_1412

//BADD_1389 replaced by BADD_1411

//BADD_1388 replaced by BADD_1410

//KaratsubaCore_701 replaced by KaratsubaCore_717

//KaratsubaCore_700 replaced by KaratsubaCore_718

//KaratsubaCore_699 replaced by KaratsubaCore_717

//BADD_1394 replaced by BADD_1406

//BADD_1393 replaced by BADD_1408

//BADD_1392 replaced by BADD_1407

//BADD_1391 replaced by BADD_1406

//KaratsubaCore_704 replaced by KaratsubaCore_718

//KaratsubaCore_703 replaced by KaratsubaCore_715

//KaratsubaCore_702 replaced by KaratsubaCore_718

//BADD_1398 replaced by BADD_1395

module BADD_1397 (
  input      [100:0]  io_a,
  input      [100:0]  io_b,
  input               io_c,
  output reg [101:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [5:0]    _zz__zz_io_s_6;
  wire       [5:0]    _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [5:0]    _zz_io_s_6;
  reg        [4:0]    _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[100 : 96]} + {1'b0,io_b[100 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {5'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[100 : 96] = _zz_io_s_7;
    io_s[101] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[4:0];
    _zz_io_s_8 <= _zz_io_s_6[5];
  end


endmodule

module BADD_1396 (
  input      [100:0]  io_a,
  input      [100:0]  io_b,
  input               io_c,
  output reg [101:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [100:0]  _zz__zz_io_s_1;
  wire       [48:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [100:0]  _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_3_3;
  wire       [0:0]    _zz__zz_io_s_3_4;
  wire       [5:0]    _zz__zz_io_s_6;
  wire       [100:0]  _zz__zz_io_s_6_1;
  wire       [5:0]    _zz__zz_io_s_6_2;
  wire       [0:0]    _zz__zz_io_s_6_3;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [5:0]    _zz_io_s_6;
  reg        [4:0]    _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,_zz__zz_io_s_1[47 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {48'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_3_1 = ({1'b0,io_a[95 : 48]} + {1'b0,_zz__zz_io_s_3_2[95 : 48]});
  assign _zz__zz_io_s_3_2 = (~ io_b);
  assign _zz__zz_io_s_3_4 = _zz_io_s_2;
  assign _zz__zz_io_s_3_3 = {48'd0, _zz__zz_io_s_3_4};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[100 : 96]} + {1'b0,_zz__zz_io_s_6_1[100 : 96]});
  assign _zz__zz_io_s_6_1 = (~ io_b);
  assign _zz__zz_io_s_6_3 = _zz_io_s_5;
  assign _zz__zz_io_s_6_2 = {5'd0, _zz__zz_io_s_6_3};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[100 : 96] = _zz_io_s_7;
    io_s[101] = (! _zz_io_s_8);
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3_1 + _zz__zz_io_s_3_3);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_2);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[4:0];
    _zz_io_s_8 <= _zz_io_s_6[5];
  end


endmodule

module BADD_1395 (
  input      [99:0]   io_a,
  input      [99:0]   io_b,
  input               io_c,
  output reg [100:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [4:0]    _zz__zz_io_s_6;
  wire       [4:0]    _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [4:0]    _zz_io_s_6;
  reg        [3:0]    _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[99 : 96]} + {1'b0,io_b[99 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {4'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[99 : 96] = _zz_io_s_7;
    io_s[100] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[3:0];
    _zz_io_s_8 <= _zz_io_s_6[4];
  end


endmodule

//KaratsubaCore_707 replaced by KaratsubaCore_715

module KaratsubaCore_706 (
  input      [50:0]   io_a_0,
  input      [50:0]   io_b_0,
  output     [101:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [101:0]  basic_mul_io_p;

  BasicMUL48_472 basic_mul (
    .io_a   (io_a_0[50:0]         ), //i
    .io_b   (io_b_0[50:0]         ), //i
    .io_p   (basic_mul_io_p[101:0]), //o
    .clk    (clk                  ), //i
    .resetn (resetn               )  //i
  );
  assign io_p = basic_mul_io_p;

endmodule

//KaratsubaCore_705 replaced by KaratsubaCore_715

//BADD_1402 replaced by BADD_1406

//BADD_1401 replaced by BADD_1408

//BADD_1400 replaced by BADD_1407

//BADD_1399 replaced by BADD_1406

//KaratsubaCore_710 replaced by KaratsubaCore_718

//KaratsubaCore_709 replaced by KaratsubaCore_715

//KaratsubaCore_708 replaced by KaratsubaCore_718

//BADD_1405 replaced by BADD_1412

//BADD_1404 replaced by BADD_1411

//BADD_1403 replaced by BADD_1410

//KaratsubaCore_713 replaced by KaratsubaCore_717

//KaratsubaCore_712 replaced by KaratsubaCore_718

//KaratsubaCore_711 replaced by KaratsubaCore_717

//BADD_1409 replaced by BADD_1406

module BADD_1408 (
  input      [98:0]   io_a,
  input      [98:0]   io_b,
  input               io_c,
  output reg [99:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [3:0]    _zz__zz_io_s_6;
  wire       [3:0]    _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [3:0]    _zz_io_s_6;
  reg        [2:0]    _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[98 : 96]} + {1'b0,io_b[98 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {3'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[98 : 96] = _zz_io_s_7;
    io_s[99] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[2:0];
    _zz_io_s_8 <= _zz_io_s_6[3];
  end


endmodule

module BADD_1407 (
  input      [98:0]   io_a,
  input      [98:0]   io_b,
  input               io_c,
  output reg [99:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [98:0]   _zz__zz_io_s_1;
  wire       [48:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [98:0]   _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_3_3;
  wire       [0:0]    _zz__zz_io_s_3_4;
  wire       [3:0]    _zz__zz_io_s_6;
  wire       [98:0]   _zz__zz_io_s_6_1;
  wire       [3:0]    _zz__zz_io_s_6_2;
  wire       [0:0]    _zz__zz_io_s_6_3;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [3:0]    _zz_io_s_6;
  reg        [2:0]    _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,_zz__zz_io_s_1[47 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {48'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_3_1 = ({1'b0,io_a[95 : 48]} + {1'b0,_zz__zz_io_s_3_2[95 : 48]});
  assign _zz__zz_io_s_3_2 = (~ io_b);
  assign _zz__zz_io_s_3_4 = _zz_io_s_2;
  assign _zz__zz_io_s_3_3 = {48'd0, _zz__zz_io_s_3_4};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[98 : 96]} + {1'b0,_zz__zz_io_s_6_1[98 : 96]});
  assign _zz__zz_io_s_6_1 = (~ io_b);
  assign _zz__zz_io_s_6_3 = _zz_io_s_5;
  assign _zz__zz_io_s_6_2 = {3'd0, _zz__zz_io_s_6_3};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[98 : 96] = _zz_io_s_7;
    io_s[99] = (! _zz_io_s_8);
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3_1 + _zz__zz_io_s_3_3);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_2);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[2:0];
    _zz_io_s_8 <= _zz_io_s_6[3];
  end


endmodule

module BADD_1406 (
  input      [97:0]   io_a,
  input      [97:0]   io_b,
  input               io_c,
  output reg [98:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [2:0]    _zz__zz_io_s_6;
  wire       [2:0]    _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [2:0]    _zz_io_s_6;
  reg        [1:0]    _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[97 : 96]} + {1'b0,io_b[97 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {2'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[97 : 96] = _zz_io_s_7;
    io_s[98] = _zz_io_s_8;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[1:0];
    _zz_io_s_8 <= _zz_io_s_6[2];
  end


endmodule

//KaratsubaCore_716 replaced by KaratsubaCore_718

module KaratsubaCore_715 (
  input      [49:0]   io_a_0,
  input      [49:0]   io_b_0,
  output     [99:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [99:0]   basic_mul_io_p;

  BasicMUL48_481 basic_mul (
    .io_a   (io_a_0[49:0]        ), //i
    .io_b   (io_b_0[49:0]        ), //i
    .io_p   (basic_mul_io_p[99:0]), //o
    .clk    (clk                 ), //i
    .resetn (resetn              )  //i
  );
  assign io_p = basic_mul_io_p;

endmodule

//KaratsubaCore_714 replaced by KaratsubaCore_718

module BADD_1412 (
  input      [143:0]  io_a,
  input      [143:0]  io_b,
  input               io_c,
  output reg [144:0]  io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_6;
  wire       [48:0]   _zz__zz_io_s_6_1;
  wire       [0:0]    _zz__zz_io_s_6_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [48:0]   _zz_io_s_6;
  reg        [47:0]   _zz_io_s_7;
  reg                 _zz_io_s_8;
  reg                 _zz_io_s_9;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[143 : 96]} + {1'b0,io_b[143 : 96]});
  assign _zz__zz_io_s_6_2 = _zz_io_s_5;
  assign _zz__zz_io_s_6_1 = {48'd0, _zz__zz_io_s_6_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[143 : 96] = _zz_io_s_7;
    io_s[144] = _zz_io_s_9;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[47:0];
    _zz_io_s_8 <= _zz_io_s_6[48];
    _zz_io_s_9 <= _zz_io_s_8;
  end


endmodule

module BADD_1411 (
  input      [96:0]   io_a,
  input      [96:0]   io_b,
  input               io_c,
  output reg [97:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [96:0]   _zz__zz_io_s_1;
  wire       [48:0]   _zz__zz_io_s_2;
  wire       [0:0]    _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [96:0]   _zz__zz_io_s_3_2;
  wire       [48:0]   _zz__zz_io_s_3_3;
  wire       [0:0]    _zz__zz_io_s_3_4;
  wire       [1:0]    _zz__zz_io_s_6;
  wire       [96:0]   _zz__zz_io_s_6_1;
  wire       [1:0]    _zz__zz_io_s_6_2;
  wire       [0:0]    _zz__zz_io_s_6_3;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  wire       [1:0]    _zz_io_s_6;
  reg        [0:0]    _zz_io_s_7;
  reg                 _zz_io_s_8;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,_zz__zz_io_s_1[47 : 0]});
  assign _zz__zz_io_s_1 = (~ io_b);
  assign _zz__zz_io_s_3 = io_c;
  assign _zz__zz_io_s_2 = {48'd0, _zz__zz_io_s_3};
  assign _zz__zz_io_s_3_1 = ({1'b0,io_a[95 : 48]} + {1'b0,_zz__zz_io_s_3_2[95 : 48]});
  assign _zz__zz_io_s_3_2 = (~ io_b);
  assign _zz__zz_io_s_3_4 = _zz_io_s_2;
  assign _zz__zz_io_s_3_3 = {48'd0, _zz__zz_io_s_3_4};
  assign _zz__zz_io_s_6 = ({1'b0,io_a[96 : 96]} + {1'b0,_zz__zz_io_s_6_1[96 : 96]});
  assign _zz__zz_io_s_6_1 = (~ io_b);
  assign _zz__zz_io_s_6_3 = _zz_io_s_5;
  assign _zz__zz_io_s_6_2 = {1'd0, _zz__zz_io_s_6_3};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_2);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[96 : 96] = _zz_io_s_7;
    io_s[97] = (! _zz_io_s_8);
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3_1 + _zz__zz_io_s_3_3);
  assign _zz_io_s_6 = (_zz__zz_io_s_6 + _zz__zz_io_s_6_2);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_7 <= _zz_io_s_6[0:0];
    _zz_io_s_8 <= _zz_io_s_6[1];
  end


endmodule

module BADD_1410 (
  input      [95:0]   io_a,
  input      [95:0]   io_b,
  input               io_c,
  output reg [96:0]   io_s,
  input               clk,
  input               resetn
);

  wire       [48:0]   _zz__zz_io_s;
  wire       [48:0]   _zz__zz_io_s_1;
  wire       [0:0]    _zz__zz_io_s_2;
  wire       [48:0]   _zz__zz_io_s_3;
  wire       [48:0]   _zz__zz_io_s_3_1;
  wire       [0:0]    _zz__zz_io_s_3_2;
  wire       [48:0]   _zz_io_s;
  reg        [47:0]   _zz_io_s_1;
  reg                 _zz_io_s_2;
  wire       [48:0]   _zz_io_s_3;
  reg        [47:0]   _zz_io_s_4;
  reg                 _zz_io_s_5;
  reg                 _zz_io_s_6;

  assign _zz__zz_io_s = ({1'b0,io_a[47 : 0]} + {1'b0,io_b[47 : 0]});
  assign _zz__zz_io_s_2 = io_c;
  assign _zz__zz_io_s_1 = {48'd0, _zz__zz_io_s_2};
  assign _zz__zz_io_s_3 = ({1'b0,io_a[95 : 48]} + {1'b0,io_b[95 : 48]});
  assign _zz__zz_io_s_3_2 = _zz_io_s_2;
  assign _zz__zz_io_s_3_1 = {48'd0, _zz__zz_io_s_3_2};
  assign _zz_io_s = (_zz__zz_io_s + _zz__zz_io_s_1);
  always @(*) begin
    io_s[47 : 0] = _zz_io_s_1;
    io_s[95 : 48] = _zz_io_s_4;
    io_s[96] = _zz_io_s_6;
  end

  assign _zz_io_s_3 = (_zz__zz_io_s_3 + _zz__zz_io_s_3_1);
  always @(posedge clk) begin
    _zz_io_s_1 <= _zz_io_s[47:0];
    _zz_io_s_2 <= _zz_io_s[48];
    _zz_io_s_4 <= _zz_io_s_3[47:0];
    _zz_io_s_5 <= _zz_io_s_3[48];
    _zz_io_s_6 <= _zz_io_s_5;
  end


endmodule

//KaratsubaCore_719 replaced by KaratsubaCore_717

module KaratsubaCore_718 (
  input      [48:0]   io_a_0,
  input      [48:0]   io_b_0,
  output     [97:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [97:0]   basic_mul_io_p;

  BasicMUL48_484 basic_mul (
    .io_a   (io_a_0[48:0]        ), //i
    .io_b   (io_b_0[48:0]        ), //i
    .io_p   (basic_mul_io_p[97:0]), //o
    .clk    (clk                 ), //i
    .resetn (resetn              )  //i
  );
  assign io_p = basic_mul_io_p;

endmodule

module KaratsubaCore_717 (
  input      [47:0]   io_a_0,
  input      [47:0]   io_b_0,
  output     [95:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [95:0]   basic_mul_io_p;

  BasicMUL48_485 basic_mul (
    .io_a   (io_a_0[47:0]        ), //i
    .io_b   (io_b_0[47:0]        ), //i
    .io_p   (basic_mul_io_p[95:0]), //o
    .clk    (clk                 ), //i
    .resetn (resetn              )  //i
  );
  assign io_p = basic_mul_io_p;

endmodule

//BasicMUL48 replaced by BasicMUL48_485

//BasicMUL48_1 replaced by BasicMUL48_484

//BasicMUL48_2 replaced by BasicMUL48_485

//BasicMUL48_3 replaced by BasicMUL48_484

//BasicMUL48_4 replaced by BasicMUL48_481

//BasicMUL48_5 replaced by BasicMUL48_484

//BasicMUL48_6 replaced by BasicMUL48_485

//BasicMUL48_7 replaced by BasicMUL48_484

//BasicMUL48_8 replaced by BasicMUL48_485

//BasicMUL48_9 replaced by BasicMUL48_484

//BasicMUL48_10 replaced by BasicMUL48_481

//BasicMUL48_11 replaced by BasicMUL48_484

//BasicMUL48_12 replaced by BasicMUL48_481

//BasicMUL48_13 replaced by BasicMUL48_472

//BasicMUL48_14 replaced by BasicMUL48_481

//BasicMUL48_15 replaced by BasicMUL48_484

//BasicMUL48_16 replaced by BasicMUL48_481

//BasicMUL48_17 replaced by BasicMUL48_484

//BasicMUL48_18 replaced by BasicMUL48_485

//BasicMUL48_19 replaced by BasicMUL48_484

//BasicMUL48_20 replaced by BasicMUL48_485

//BasicMUL48_21 replaced by BasicMUL48_484

//BasicMUL48_22 replaced by BasicMUL48_481

//BasicMUL48_23 replaced by BasicMUL48_484

//BasicMUL48_24 replaced by BasicMUL48_485

//BasicMUL48_25 replaced by BasicMUL48_484

//BasicMUL48_26 replaced by BasicMUL48_485

//BasicMUL48_27 replaced by BasicMUL48_485

//BasicMUL48_28 replaced by BasicMUL48_484

//BasicMUL48_29 replaced by BasicMUL48_485

//BasicMUL48_30 replaced by BasicMUL48_484

//BasicMUL48_31 replaced by BasicMUL48_481

//BasicMUL48_32 replaced by BasicMUL48_484

//BasicMUL48_33 replaced by BasicMUL48_485

//BasicMUL48_34 replaced by BasicMUL48_484

//BasicMUL48_35 replaced by BasicMUL48_485

//BasicMUL48_36 replaced by BasicMUL48_484

//BasicMUL48_37 replaced by BasicMUL48_481

//BasicMUL48_38 replaced by BasicMUL48_484

//BasicMUL48_39 replaced by BasicMUL48_481

//BasicMUL48_40 replaced by BasicMUL48_472

//BasicMUL48_41 replaced by BasicMUL48_481

//BasicMUL48_42 replaced by BasicMUL48_484

//BasicMUL48_43 replaced by BasicMUL48_481

//BasicMUL48_44 replaced by BasicMUL48_484

//BasicMUL48_45 replaced by BasicMUL48_485

//BasicMUL48_46 replaced by BasicMUL48_484

//BasicMUL48_47 replaced by BasicMUL48_485

//BasicMUL48_48 replaced by BasicMUL48_484

//BasicMUL48_49 replaced by BasicMUL48_481

//BasicMUL48_50 replaced by BasicMUL48_484

//BasicMUL48_51 replaced by BasicMUL48_485

//BasicMUL48_52 replaced by BasicMUL48_484

//BasicMUL48_53 replaced by BasicMUL48_485

//BasicMUL48_54 replaced by BasicMUL48_485

//BasicMUL48_55 replaced by BasicMUL48_484

//BasicMUL48_56 replaced by BasicMUL48_485

//BasicMUL48_57 replaced by BasicMUL48_484

//BasicMUL48_58 replaced by BasicMUL48_481

//BasicMUL48_59 replaced by BasicMUL48_484

//BasicMUL48_60 replaced by BasicMUL48_485

//BasicMUL48_61 replaced by BasicMUL48_484

//BasicMUL48_62 replaced by BasicMUL48_485

//BasicMUL48_63 replaced by BasicMUL48_484

//BasicMUL48_64 replaced by BasicMUL48_481

//BasicMUL48_65 replaced by BasicMUL48_484

//BasicMUL48_66 replaced by BasicMUL48_481

//BasicMUL48_67 replaced by BasicMUL48_472

//BasicMUL48_68 replaced by BasicMUL48_481

//BasicMUL48_69 replaced by BasicMUL48_484

//BasicMUL48_70 replaced by BasicMUL48_481

//BasicMUL48_71 replaced by BasicMUL48_484

//BasicMUL48_72 replaced by BasicMUL48_485

//BasicMUL48_73 replaced by BasicMUL48_484

//BasicMUL48_74 replaced by BasicMUL48_485

//BasicMUL48_75 replaced by BasicMUL48_484

//BasicMUL48_76 replaced by BasicMUL48_481

//BasicMUL48_77 replaced by BasicMUL48_484

//BasicMUL48_78 replaced by BasicMUL48_485

//BasicMUL48_79 replaced by BasicMUL48_484

//BasicMUL48_80 replaced by BasicMUL48_485

//BasicMUL48_81 replaced by BasicMUL48_485

//BasicMUL48_82 replaced by BasicMUL48_484

//BasicMUL48_83 replaced by BasicMUL48_485

//BasicMUL48_84 replaced by BasicMUL48_484

//BasicMUL48_85 replaced by BasicMUL48_481

//BasicMUL48_86 replaced by BasicMUL48_484

//BasicMUL48_87 replaced by BasicMUL48_485

//BasicMUL48_88 replaced by BasicMUL48_484

//BasicMUL48_89 replaced by BasicMUL48_485

//BasicMUL48_90 replaced by BasicMUL48_484

//BasicMUL48_91 replaced by BasicMUL48_481

//BasicMUL48_92 replaced by BasicMUL48_484

//BasicMUL48_93 replaced by BasicMUL48_481

//BasicMUL48_94 replaced by BasicMUL48_472

//BasicMUL48_95 replaced by BasicMUL48_481

//BasicMUL48_96 replaced by BasicMUL48_484

//BasicMUL48_97 replaced by BasicMUL48_481

//BasicMUL48_98 replaced by BasicMUL48_484

//BasicMUL48_99 replaced by BasicMUL48_485

//BasicMUL48_100 replaced by BasicMUL48_484

//BasicMUL48_101 replaced by BasicMUL48_485

//BasicMUL48_102 replaced by BasicMUL48_484

//BasicMUL48_103 replaced by BasicMUL48_481

//BasicMUL48_104 replaced by BasicMUL48_484

//BasicMUL48_105 replaced by BasicMUL48_485

//BasicMUL48_106 replaced by BasicMUL48_484

//BasicMUL48_107 replaced by BasicMUL48_485

//BasicMUL48_108 replaced by BasicMUL48_485

//BasicMUL48_109 replaced by BasicMUL48_484

//BasicMUL48_110 replaced by BasicMUL48_485

//BasicMUL48_111 replaced by BasicMUL48_484

//BasicMUL48_112 replaced by BasicMUL48_481

//BasicMUL48_113 replaced by BasicMUL48_484

//BasicMUL48_114 replaced by BasicMUL48_485

//BasicMUL48_115 replaced by BasicMUL48_484

//BasicMUL48_116 replaced by BasicMUL48_485

//BasicMUL48_117 replaced by BasicMUL48_484

//BasicMUL48_118 replaced by BasicMUL48_481

//BasicMUL48_119 replaced by BasicMUL48_484

//BasicMUL48_120 replaced by BasicMUL48_481

//BasicMUL48_121 replaced by BasicMUL48_472

//BasicMUL48_122 replaced by BasicMUL48_481

//BasicMUL48_123 replaced by BasicMUL48_484

//BasicMUL48_124 replaced by BasicMUL48_481

//BasicMUL48_125 replaced by BasicMUL48_484

//BasicMUL48_126 replaced by BasicMUL48_485

//BasicMUL48_127 replaced by BasicMUL48_484

//BasicMUL48_128 replaced by BasicMUL48_485

//BasicMUL48_129 replaced by BasicMUL48_484

//BasicMUL48_130 replaced by BasicMUL48_481

//BasicMUL48_131 replaced by BasicMUL48_484

//BasicMUL48_132 replaced by BasicMUL48_485

//BasicMUL48_133 replaced by BasicMUL48_484

//BasicMUL48_134 replaced by BasicMUL48_485

//BasicMUL48_135 replaced by BasicMUL48_485

//BasicMUL48_136 replaced by BasicMUL48_484

//BasicMUL48_137 replaced by BasicMUL48_485

//BasicMUL48_138 replaced by BasicMUL48_484

//BasicMUL48_139 replaced by BasicMUL48_481

//BasicMUL48_140 replaced by BasicMUL48_484

//BasicMUL48_141 replaced by BasicMUL48_485

//BasicMUL48_142 replaced by BasicMUL48_484

//BasicMUL48_143 replaced by BasicMUL48_485

//BasicMUL48_144 replaced by BasicMUL48_484

//BasicMUL48_145 replaced by BasicMUL48_481

//BasicMUL48_146 replaced by BasicMUL48_484

//BasicMUL48_147 replaced by BasicMUL48_481

//BasicMUL48_148 replaced by BasicMUL48_472

//BasicMUL48_149 replaced by BasicMUL48_481

//BasicMUL48_150 replaced by BasicMUL48_484

//BasicMUL48_151 replaced by BasicMUL48_481

//BasicMUL48_152 replaced by BasicMUL48_484

//BasicMUL48_153 replaced by BasicMUL48_485

//BasicMUL48_154 replaced by BasicMUL48_484

//BasicMUL48_155 replaced by BasicMUL48_485

//BasicMUL48_156 replaced by BasicMUL48_484

//BasicMUL48_157 replaced by BasicMUL48_481

//BasicMUL48_158 replaced by BasicMUL48_484

//BasicMUL48_159 replaced by BasicMUL48_485

//BasicMUL48_160 replaced by BasicMUL48_484

//BasicMUL48_161 replaced by BasicMUL48_485

//BasicMUL48_162 replaced by BasicMUL48_485

//BasicMUL48_163 replaced by BasicMUL48_484

//BasicMUL48_164 replaced by BasicMUL48_485

//BasicMUL48_165 replaced by BasicMUL48_484

//BasicMUL48_166 replaced by BasicMUL48_481

//BasicMUL48_167 replaced by BasicMUL48_484

//BasicMUL48_168 replaced by BasicMUL48_485

//BasicMUL48_169 replaced by BasicMUL48_484

//BasicMUL48_170 replaced by BasicMUL48_485

//BasicMUL48_171 replaced by BasicMUL48_484

//BasicMUL48_172 replaced by BasicMUL48_481

//BasicMUL48_173 replaced by BasicMUL48_484

//BasicMUL48_174 replaced by BasicMUL48_481

//BasicMUL48_175 replaced by BasicMUL48_472

//BasicMUL48_176 replaced by BasicMUL48_481

//BasicMUL48_177 replaced by BasicMUL48_484

//BasicMUL48_178 replaced by BasicMUL48_481

//BasicMUL48_179 replaced by BasicMUL48_484

//BasicMUL48_180 replaced by BasicMUL48_485

//BasicMUL48_181 replaced by BasicMUL48_484

//BasicMUL48_182 replaced by BasicMUL48_485

//BasicMUL48_183 replaced by BasicMUL48_484

//BasicMUL48_184 replaced by BasicMUL48_481

//BasicMUL48_185 replaced by BasicMUL48_484

//BasicMUL48_186 replaced by BasicMUL48_485

//BasicMUL48_187 replaced by BasicMUL48_484

//BasicMUL48_188 replaced by BasicMUL48_485

//BasicMUL48_189 replaced by BasicMUL48_485

//BasicMUL48_190 replaced by BasicMUL48_484

//BasicMUL48_191 replaced by BasicMUL48_485

//BasicMUL48_192 replaced by BasicMUL48_484

//BasicMUL48_193 replaced by BasicMUL48_481

//BasicMUL48_194 replaced by BasicMUL48_484

//BasicMUL48_195 replaced by BasicMUL48_485

//BasicMUL48_196 replaced by BasicMUL48_484

//BasicMUL48_197 replaced by BasicMUL48_485

//BasicMUL48_198 replaced by BasicMUL48_484

//BasicMUL48_199 replaced by BasicMUL48_481

//BasicMUL48_200 replaced by BasicMUL48_484

//BasicMUL48_201 replaced by BasicMUL48_481

//BasicMUL48_202 replaced by BasicMUL48_472

//BasicMUL48_203 replaced by BasicMUL48_481

//BasicMUL48_204 replaced by BasicMUL48_484

//BasicMUL48_205 replaced by BasicMUL48_481

//BasicMUL48_206 replaced by BasicMUL48_484

//BasicMUL48_207 replaced by BasicMUL48_485

//BasicMUL48_208 replaced by BasicMUL48_484

//BasicMUL48_209 replaced by BasicMUL48_485

//BasicMUL48_210 replaced by BasicMUL48_484

//BasicMUL48_211 replaced by BasicMUL48_481

//BasicMUL48_212 replaced by BasicMUL48_484

//BasicMUL48_213 replaced by BasicMUL48_485

//BasicMUL48_214 replaced by BasicMUL48_484

//BasicMUL48_215 replaced by BasicMUL48_485

//BasicMUL48_216 replaced by BasicMUL48_485

//BasicMUL48_217 replaced by BasicMUL48_484

//BasicMUL48_218 replaced by BasicMUL48_485

//BasicMUL48_219 replaced by BasicMUL48_484

//BasicMUL48_220 replaced by BasicMUL48_481

//BasicMUL48_221 replaced by BasicMUL48_484

//BasicMUL48_222 replaced by BasicMUL48_485

//BasicMUL48_223 replaced by BasicMUL48_484

//BasicMUL48_224 replaced by BasicMUL48_485

//BasicMUL48_225 replaced by BasicMUL48_484

//BasicMUL48_226 replaced by BasicMUL48_481

//BasicMUL48_227 replaced by BasicMUL48_484

//BasicMUL48_228 replaced by BasicMUL48_481

//BasicMUL48_229 replaced by BasicMUL48_472

//BasicMUL48_230 replaced by BasicMUL48_481

//BasicMUL48_231 replaced by BasicMUL48_484

//BasicMUL48_232 replaced by BasicMUL48_481

//BasicMUL48_233 replaced by BasicMUL48_484

//BasicMUL48_234 replaced by BasicMUL48_485

//BasicMUL48_235 replaced by BasicMUL48_484

//BasicMUL48_236 replaced by BasicMUL48_485

//BasicMUL48_237 replaced by BasicMUL48_484

//BasicMUL48_238 replaced by BasicMUL48_481

//BasicMUL48_239 replaced by BasicMUL48_484

//BasicMUL48_240 replaced by BasicMUL48_485

//BasicMUL48_241 replaced by BasicMUL48_484

//BasicMUL48_242 replaced by BasicMUL48_485

//BasicMUL48_243 replaced by BasicMUL48_485

//BasicMUL48_244 replaced by BasicMUL48_484

//BasicMUL48_245 replaced by BasicMUL48_485

//BasicMUL48_246 replaced by BasicMUL48_484

//BasicMUL48_247 replaced by BasicMUL48_481

//BasicMUL48_248 replaced by BasicMUL48_484

//BasicMUL48_249 replaced by BasicMUL48_485

//BasicMUL48_250 replaced by BasicMUL48_484

//BasicMUL48_251 replaced by BasicMUL48_485

//BasicMUL48_252 replaced by BasicMUL48_484

//BasicMUL48_253 replaced by BasicMUL48_481

//BasicMUL48_254 replaced by BasicMUL48_484

//BasicMUL48_255 replaced by BasicMUL48_481

//BasicMUL48_256 replaced by BasicMUL48_472

//BasicMUL48_257 replaced by BasicMUL48_481

//BasicMUL48_258 replaced by BasicMUL48_484

//BasicMUL48_259 replaced by BasicMUL48_481

//BasicMUL48_260 replaced by BasicMUL48_484

//BasicMUL48_261 replaced by BasicMUL48_485

//BasicMUL48_262 replaced by BasicMUL48_484

//BasicMUL48_263 replaced by BasicMUL48_485

//BasicMUL48_264 replaced by BasicMUL48_484

//BasicMUL48_265 replaced by BasicMUL48_481

//BasicMUL48_266 replaced by BasicMUL48_484

//BasicMUL48_267 replaced by BasicMUL48_485

//BasicMUL48_268 replaced by BasicMUL48_484

//BasicMUL48_269 replaced by BasicMUL48_485

//BasicMUL48_270 replaced by BasicMUL48_485

//BasicMUL48_271 replaced by BasicMUL48_484

//BasicMUL48_272 replaced by BasicMUL48_485

//BasicMUL48_273 replaced by BasicMUL48_484

//BasicMUL48_274 replaced by BasicMUL48_481

//BasicMUL48_275 replaced by BasicMUL48_484

//BasicMUL48_276 replaced by BasicMUL48_485

//BasicMUL48_277 replaced by BasicMUL48_484

//BasicMUL48_278 replaced by BasicMUL48_485

//BasicMUL48_279 replaced by BasicMUL48_484

//BasicMUL48_280 replaced by BasicMUL48_481

//BasicMUL48_281 replaced by BasicMUL48_484

//BasicMUL48_282 replaced by BasicMUL48_481

//BasicMUL48_283 replaced by BasicMUL48_472

//BasicMUL48_284 replaced by BasicMUL48_481

//BasicMUL48_285 replaced by BasicMUL48_484

//BasicMUL48_286 replaced by BasicMUL48_481

//BasicMUL48_287 replaced by BasicMUL48_484

//BasicMUL48_288 replaced by BasicMUL48_485

//BasicMUL48_289 replaced by BasicMUL48_484

//BasicMUL48_290 replaced by BasicMUL48_485

//BasicMUL48_291 replaced by BasicMUL48_484

//BasicMUL48_292 replaced by BasicMUL48_481

//BasicMUL48_293 replaced by BasicMUL48_484

//BasicMUL48_294 replaced by BasicMUL48_485

//BasicMUL48_295 replaced by BasicMUL48_484

//BasicMUL48_296 replaced by BasicMUL48_485

//BasicMUL48_297 replaced by BasicMUL48_485

//BasicMUL48_298 replaced by BasicMUL48_484

//BasicMUL48_299 replaced by BasicMUL48_485

//BasicMUL48_300 replaced by BasicMUL48_484

//BasicMUL48_301 replaced by BasicMUL48_481

//BasicMUL48_302 replaced by BasicMUL48_484

//BasicMUL48_303 replaced by BasicMUL48_485

//BasicMUL48_304 replaced by BasicMUL48_484

//BasicMUL48_305 replaced by BasicMUL48_485

//BasicMUL48_306 replaced by BasicMUL48_484

//BasicMUL48_307 replaced by BasicMUL48_481

//BasicMUL48_308 replaced by BasicMUL48_484

//BasicMUL48_309 replaced by BasicMUL48_481

//BasicMUL48_310 replaced by BasicMUL48_472

//BasicMUL48_311 replaced by BasicMUL48_481

//BasicMUL48_312 replaced by BasicMUL48_484

//BasicMUL48_313 replaced by BasicMUL48_481

//BasicMUL48_314 replaced by BasicMUL48_484

//BasicMUL48_315 replaced by BasicMUL48_485

//BasicMUL48_316 replaced by BasicMUL48_484

//BasicMUL48_317 replaced by BasicMUL48_485

//BasicMUL48_318 replaced by BasicMUL48_484

//BasicMUL48_319 replaced by BasicMUL48_481

//BasicMUL48_320 replaced by BasicMUL48_484

//BasicMUL48_321 replaced by BasicMUL48_485

//BasicMUL48_322 replaced by BasicMUL48_484

//BasicMUL48_323 replaced by BasicMUL48_485

//BasicMUL48_324 replaced by BasicMUL48_485

//BasicMUL48_325 replaced by BasicMUL48_484

//BasicMUL48_326 replaced by BasicMUL48_485

//BasicMUL48_327 replaced by BasicMUL48_484

//BasicMUL48_328 replaced by BasicMUL48_481

//BasicMUL48_329 replaced by BasicMUL48_484

//BasicMUL48_330 replaced by BasicMUL48_485

//BasicMUL48_331 replaced by BasicMUL48_484

//BasicMUL48_332 replaced by BasicMUL48_485

//BasicMUL48_333 replaced by BasicMUL48_484

//BasicMUL48_334 replaced by BasicMUL48_481

//BasicMUL48_335 replaced by BasicMUL48_484

//BasicMUL48_336 replaced by BasicMUL48_481

//BasicMUL48_337 replaced by BasicMUL48_472

//BasicMUL48_338 replaced by BasicMUL48_481

//BasicMUL48_339 replaced by BasicMUL48_484

//BasicMUL48_340 replaced by BasicMUL48_481

//BasicMUL48_341 replaced by BasicMUL48_484

//BasicMUL48_342 replaced by BasicMUL48_485

//BasicMUL48_343 replaced by BasicMUL48_484

//BasicMUL48_344 replaced by BasicMUL48_485

//BasicMUL48_345 replaced by BasicMUL48_484

//BasicMUL48_346 replaced by BasicMUL48_481

//BasicMUL48_347 replaced by BasicMUL48_484

//BasicMUL48_348 replaced by BasicMUL48_485

//BasicMUL48_349 replaced by BasicMUL48_484

//BasicMUL48_350 replaced by BasicMUL48_485

//BasicMUL48_351 replaced by BasicMUL48_485

//BasicMUL48_352 replaced by BasicMUL48_484

//BasicMUL48_353 replaced by BasicMUL48_485

//BasicMUL48_354 replaced by BasicMUL48_484

//BasicMUL48_355 replaced by BasicMUL48_481

//BasicMUL48_356 replaced by BasicMUL48_484

//BasicMUL48_357 replaced by BasicMUL48_485

//BasicMUL48_358 replaced by BasicMUL48_484

//BasicMUL48_359 replaced by BasicMUL48_485

//BasicMUL48_360 replaced by BasicMUL48_484

//BasicMUL48_361 replaced by BasicMUL48_481

//BasicMUL48_362 replaced by BasicMUL48_484

//BasicMUL48_363 replaced by BasicMUL48_481

//BasicMUL48_364 replaced by BasicMUL48_472

//BasicMUL48_365 replaced by BasicMUL48_481

//BasicMUL48_366 replaced by BasicMUL48_484

//BasicMUL48_367 replaced by BasicMUL48_481

//BasicMUL48_368 replaced by BasicMUL48_484

//BasicMUL48_369 replaced by BasicMUL48_485

//BasicMUL48_370 replaced by BasicMUL48_484

//BasicMUL48_371 replaced by BasicMUL48_485

//BasicMUL48_372 replaced by BasicMUL48_484

//BasicMUL48_373 replaced by BasicMUL48_481

//BasicMUL48_374 replaced by BasicMUL48_484

//BasicMUL48_375 replaced by BasicMUL48_485

//BasicMUL48_376 replaced by BasicMUL48_484

//BasicMUL48_377 replaced by BasicMUL48_485

//BasicMUL48_378 replaced by BasicMUL48_485

//BasicMUL48_379 replaced by BasicMUL48_484

//BasicMUL48_380 replaced by BasicMUL48_485

//BasicMUL48_381 replaced by BasicMUL48_484

//BasicMUL48_382 replaced by BasicMUL48_481

//BasicMUL48_383 replaced by BasicMUL48_484

//BasicMUL48_384 replaced by BasicMUL48_485

//BasicMUL48_385 replaced by BasicMUL48_484

//BasicMUL48_386 replaced by BasicMUL48_485

//BasicMUL48_387 replaced by BasicMUL48_484

//BasicMUL48_388 replaced by BasicMUL48_481

//BasicMUL48_389 replaced by BasicMUL48_484

//BasicMUL48_390 replaced by BasicMUL48_481

//BasicMUL48_391 replaced by BasicMUL48_472

//BasicMUL48_392 replaced by BasicMUL48_481

//BasicMUL48_393 replaced by BasicMUL48_484

//BasicMUL48_394 replaced by BasicMUL48_481

//BasicMUL48_395 replaced by BasicMUL48_484

//BasicMUL48_396 replaced by BasicMUL48_485

//BasicMUL48_397 replaced by BasicMUL48_484

//BasicMUL48_398 replaced by BasicMUL48_485

//BasicMUL48_399 replaced by BasicMUL48_484

//BasicMUL48_400 replaced by BasicMUL48_481

//BasicMUL48_401 replaced by BasicMUL48_484

//BasicMUL48_402 replaced by BasicMUL48_485

//BasicMUL48_403 replaced by BasicMUL48_484

//BasicMUL48_404 replaced by BasicMUL48_485

//BasicMUL48_405 replaced by BasicMUL48_485

//BasicMUL48_406 replaced by BasicMUL48_484

//BasicMUL48_407 replaced by BasicMUL48_485

//BasicMUL48_408 replaced by BasicMUL48_484

//BasicMUL48_409 replaced by BasicMUL48_481

//BasicMUL48_410 replaced by BasicMUL48_484

//BasicMUL48_411 replaced by BasicMUL48_485

//BasicMUL48_412 replaced by BasicMUL48_484

//BasicMUL48_413 replaced by BasicMUL48_485

//BasicMUL48_414 replaced by BasicMUL48_484

//BasicMUL48_415 replaced by BasicMUL48_481

//BasicMUL48_416 replaced by BasicMUL48_484

//BasicMUL48_417 replaced by BasicMUL48_481

//BasicMUL48_418 replaced by BasicMUL48_472

//BasicMUL48_419 replaced by BasicMUL48_481

//BasicMUL48_420 replaced by BasicMUL48_484

//BasicMUL48_421 replaced by BasicMUL48_481

//BasicMUL48_422 replaced by BasicMUL48_484

//BasicMUL48_423 replaced by BasicMUL48_485

//BasicMUL48_424 replaced by BasicMUL48_484

//BasicMUL48_425 replaced by BasicMUL48_485

//BasicMUL48_426 replaced by BasicMUL48_484

//BasicMUL48_427 replaced by BasicMUL48_481

//BasicMUL48_428 replaced by BasicMUL48_484

//BasicMUL48_429 replaced by BasicMUL48_485

//BasicMUL48_430 replaced by BasicMUL48_484

//BasicMUL48_431 replaced by BasicMUL48_485

//BasicMUL48_432 replaced by BasicMUL48_485

//BasicMUL48_433 replaced by BasicMUL48_484

//BasicMUL48_434 replaced by BasicMUL48_485

//BasicMUL48_435 replaced by BasicMUL48_484

//BasicMUL48_436 replaced by BasicMUL48_481

//BasicMUL48_437 replaced by BasicMUL48_484

//BasicMUL48_438 replaced by BasicMUL48_485

//BasicMUL48_439 replaced by BasicMUL48_484

//BasicMUL48_440 replaced by BasicMUL48_485

//BasicMUL48_441 replaced by BasicMUL48_484

//BasicMUL48_442 replaced by BasicMUL48_481

//BasicMUL48_443 replaced by BasicMUL48_484

//BasicMUL48_444 replaced by BasicMUL48_481

//BasicMUL48_445 replaced by BasicMUL48_472

//BasicMUL48_446 replaced by BasicMUL48_481

//BasicMUL48_447 replaced by BasicMUL48_484

//BasicMUL48_448 replaced by BasicMUL48_481

//BasicMUL48_449 replaced by BasicMUL48_484

//BasicMUL48_450 replaced by BasicMUL48_485

//BasicMUL48_451 replaced by BasicMUL48_484

//BasicMUL48_452 replaced by BasicMUL48_485

//BasicMUL48_453 replaced by BasicMUL48_484

//BasicMUL48_454 replaced by BasicMUL48_481

//BasicMUL48_455 replaced by BasicMUL48_484

//BasicMUL48_456 replaced by BasicMUL48_485

//BasicMUL48_457 replaced by BasicMUL48_484

//BasicMUL48_458 replaced by BasicMUL48_485

//BasicMUL48_459 replaced by BasicMUL48_485

//BasicMUL48_460 replaced by BasicMUL48_484

//BasicMUL48_461 replaced by BasicMUL48_485

//BasicMUL48_462 replaced by BasicMUL48_484

//BasicMUL48_463 replaced by BasicMUL48_481

//BasicMUL48_464 replaced by BasicMUL48_484

//BasicMUL48_465 replaced by BasicMUL48_485

//BasicMUL48_466 replaced by BasicMUL48_484

//BasicMUL48_467 replaced by BasicMUL48_485

//BasicMUL48_468 replaced by BasicMUL48_484

//BasicMUL48_469 replaced by BasicMUL48_481

//BasicMUL48_470 replaced by BasicMUL48_484

//BasicMUL48_471 replaced by BasicMUL48_481

module BasicMUL48_472 (
  input      [50:0]   io_a,
  input      [50:0]   io_b,
  output     [101:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [51:0]   mul_io_a;
  wire       [102:0]  mul_io_p;
  wire       [101:0]  p;

  BasicMAC48_485 mul (
    .io_a   (mul_io_a[51:0] ), //i
    .io_b   (io_b[50:0]     ), //i
    .io_c   (51'h0          ), //i
    .io_ce  (1'b1           ), //i
    .io_p   (mul_io_p[102:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  assign io_p = p;
  assign mul_io_a = {1'd0, io_a};
  assign p = mul_io_p[101:0];

endmodule

//BasicMUL48_473 replaced by BasicMUL48_481

//BasicMUL48_474 replaced by BasicMUL48_484

//BasicMUL48_475 replaced by BasicMUL48_481

//BasicMUL48_476 replaced by BasicMUL48_484

//BasicMUL48_477 replaced by BasicMUL48_485

//BasicMUL48_478 replaced by BasicMUL48_484

//BasicMUL48_479 replaced by BasicMUL48_485

//BasicMUL48_480 replaced by BasicMUL48_484

module BasicMUL48_481 (
  input      [49:0]   io_a,
  input      [49:0]   io_b,
  output     [99:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [51:0]   mul_io_a;
  wire       [50:0]   mul_io_b;
  wire       [102:0]  mul_io_p;
  wire       [99:0]   p;

  BasicMAC48_485 mul (
    .io_a   (mul_io_a[51:0] ), //i
    .io_b   (mul_io_b[50:0] ), //i
    .io_c   (51'h0          ), //i
    .io_ce  (1'b1           ), //i
    .io_p   (mul_io_p[102:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  assign io_p = p;
  assign mul_io_a = {2'd0, io_a};
  assign mul_io_b = {1'd0, io_b};
  assign p = mul_io_p[99:0];

endmodule

//BasicMUL48_482 replaced by BasicMUL48_484

//BasicMUL48_483 replaced by BasicMUL48_485

module BasicMUL48_484 (
  input      [48:0]   io_a,
  input      [48:0]   io_b,
  output     [97:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [51:0]   mul_io_a;
  wire       [50:0]   mul_io_b;
  wire       [102:0]  mul_io_p;
  wire       [97:0]   p;

  BasicMAC48_485 mul (
    .io_a   (mul_io_a[51:0] ), //i
    .io_b   (mul_io_b[50:0] ), //i
    .io_c   (51'h0          ), //i
    .io_ce  (1'b1           ), //i
    .io_p   (mul_io_p[102:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  assign io_p = p;
  assign mul_io_a = {3'd0, io_a};
  assign mul_io_b = {2'd0, io_b};
  assign p = mul_io_p[97:0];

endmodule

module BasicMUL48_485 (
  input      [47:0]   io_a,
  input      [47:0]   io_b,
  output     [95:0]   io_p,
  input               clk,
  input               resetn
);

  wire       [51:0]   mul_io_a;
  wire       [50:0]   mul_io_b;
  wire       [102:0]  mul_io_p;
  wire       [95:0]   p;

  BasicMAC48_485 mul (
    .io_a   (mul_io_a[51:0] ), //i
    .io_b   (mul_io_b[50:0] ), //i
    .io_c   (51'h0          ), //i
    .io_ce  (1'b1           ), //i
    .io_p   (mul_io_p[102:0]), //o
    .clk    (clk            ), //i
    .resetn (resetn         )  //i
  );
  assign io_p = p;
  assign mul_io_a = {4'd0, io_a};
  assign mul_io_b = {3'd0, io_b};
  assign p = mul_io_p[95:0];

endmodule

//BasicMAC48 replaced by BasicMAC48_485

//BasicMAC48_1 replaced by BasicMAC48_485

//BasicMAC48_2 replaced by BasicMAC48_485

//BasicMAC48_3 replaced by BasicMAC48_485

//BasicMAC48_4 replaced by BasicMAC48_485

//BasicMAC48_5 replaced by BasicMAC48_485

//BasicMAC48_6 replaced by BasicMAC48_485

//BasicMAC48_7 replaced by BasicMAC48_485

//BasicMAC48_8 replaced by BasicMAC48_485

//BasicMAC48_9 replaced by BasicMAC48_485

//BasicMAC48_10 replaced by BasicMAC48_485

//BasicMAC48_11 replaced by BasicMAC48_485

//BasicMAC48_12 replaced by BasicMAC48_485

//BasicMAC48_13 replaced by BasicMAC48_485

//BasicMAC48_14 replaced by BasicMAC48_485

//BasicMAC48_15 replaced by BasicMAC48_485

//BasicMAC48_16 replaced by BasicMAC48_485

//BasicMAC48_17 replaced by BasicMAC48_485

//BasicMAC48_18 replaced by BasicMAC48_485

//BasicMAC48_19 replaced by BasicMAC48_485

//BasicMAC48_20 replaced by BasicMAC48_485

//BasicMAC48_21 replaced by BasicMAC48_485

//BasicMAC48_22 replaced by BasicMAC48_485

//BasicMAC48_23 replaced by BasicMAC48_485

//BasicMAC48_24 replaced by BasicMAC48_485

//BasicMAC48_25 replaced by BasicMAC48_485

//BasicMAC48_26 replaced by BasicMAC48_485

//BasicMAC48_27 replaced by BasicMAC48_485

//BasicMAC48_28 replaced by BasicMAC48_485

//BasicMAC48_29 replaced by BasicMAC48_485

//BasicMAC48_30 replaced by BasicMAC48_485

//BasicMAC48_31 replaced by BasicMAC48_485

//BasicMAC48_32 replaced by BasicMAC48_485

//BasicMAC48_33 replaced by BasicMAC48_485

//BasicMAC48_34 replaced by BasicMAC48_485

//BasicMAC48_35 replaced by BasicMAC48_485

//BasicMAC48_36 replaced by BasicMAC48_485

//BasicMAC48_37 replaced by BasicMAC48_485

//BasicMAC48_38 replaced by BasicMAC48_485

//BasicMAC48_39 replaced by BasicMAC48_485

//BasicMAC48_40 replaced by BasicMAC48_485

//BasicMAC48_41 replaced by BasicMAC48_485

//BasicMAC48_42 replaced by BasicMAC48_485

//BasicMAC48_43 replaced by BasicMAC48_485

//BasicMAC48_44 replaced by BasicMAC48_485

//BasicMAC48_45 replaced by BasicMAC48_485

//BasicMAC48_46 replaced by BasicMAC48_485

//BasicMAC48_47 replaced by BasicMAC48_485

//BasicMAC48_48 replaced by BasicMAC48_485

//BasicMAC48_49 replaced by BasicMAC48_485

//BasicMAC48_50 replaced by BasicMAC48_485

//BasicMAC48_51 replaced by BasicMAC48_485

//BasicMAC48_52 replaced by BasicMAC48_485

//BasicMAC48_53 replaced by BasicMAC48_485

//BasicMAC48_54 replaced by BasicMAC48_485

//BasicMAC48_55 replaced by BasicMAC48_485

//BasicMAC48_56 replaced by BasicMAC48_485

//BasicMAC48_57 replaced by BasicMAC48_485

//BasicMAC48_58 replaced by BasicMAC48_485

//BasicMAC48_59 replaced by BasicMAC48_485

//BasicMAC48_60 replaced by BasicMAC48_485

//BasicMAC48_61 replaced by BasicMAC48_485

//BasicMAC48_62 replaced by BasicMAC48_485

//BasicMAC48_63 replaced by BasicMAC48_485

//BasicMAC48_64 replaced by BasicMAC48_485

//BasicMAC48_65 replaced by BasicMAC48_485

//BasicMAC48_66 replaced by BasicMAC48_485

//BasicMAC48_67 replaced by BasicMAC48_485

//BasicMAC48_68 replaced by BasicMAC48_485

//BasicMAC48_69 replaced by BasicMAC48_485

//BasicMAC48_70 replaced by BasicMAC48_485

//BasicMAC48_71 replaced by BasicMAC48_485

//BasicMAC48_72 replaced by BasicMAC48_485

//BasicMAC48_73 replaced by BasicMAC48_485

//BasicMAC48_74 replaced by BasicMAC48_485

//BasicMAC48_75 replaced by BasicMAC48_485

//BasicMAC48_76 replaced by BasicMAC48_485

//BasicMAC48_77 replaced by BasicMAC48_485

//BasicMAC48_78 replaced by BasicMAC48_485

//BasicMAC48_79 replaced by BasicMAC48_485

//BasicMAC48_80 replaced by BasicMAC48_485

//BasicMAC48_81 replaced by BasicMAC48_485

//BasicMAC48_82 replaced by BasicMAC48_485

//BasicMAC48_83 replaced by BasicMAC48_485

//BasicMAC48_84 replaced by BasicMAC48_485

//BasicMAC48_85 replaced by BasicMAC48_485

//BasicMAC48_86 replaced by BasicMAC48_485

//BasicMAC48_87 replaced by BasicMAC48_485

//BasicMAC48_88 replaced by BasicMAC48_485

//BasicMAC48_89 replaced by BasicMAC48_485

//BasicMAC48_90 replaced by BasicMAC48_485

//BasicMAC48_91 replaced by BasicMAC48_485

//BasicMAC48_92 replaced by BasicMAC48_485

//BasicMAC48_93 replaced by BasicMAC48_485

//BasicMAC48_94 replaced by BasicMAC48_485

//BasicMAC48_95 replaced by BasicMAC48_485

//BasicMAC48_96 replaced by BasicMAC48_485

//BasicMAC48_97 replaced by BasicMAC48_485

//BasicMAC48_98 replaced by BasicMAC48_485

//BasicMAC48_99 replaced by BasicMAC48_485

//BasicMAC48_100 replaced by BasicMAC48_485

//BasicMAC48_101 replaced by BasicMAC48_485

//BasicMAC48_102 replaced by BasicMAC48_485

//BasicMAC48_103 replaced by BasicMAC48_485

//BasicMAC48_104 replaced by BasicMAC48_485

//BasicMAC48_105 replaced by BasicMAC48_485

//BasicMAC48_106 replaced by BasicMAC48_485

//BasicMAC48_107 replaced by BasicMAC48_485

//BasicMAC48_108 replaced by BasicMAC48_485

//BasicMAC48_109 replaced by BasicMAC48_485

//BasicMAC48_110 replaced by BasicMAC48_485

//BasicMAC48_111 replaced by BasicMAC48_485

//BasicMAC48_112 replaced by BasicMAC48_485

//BasicMAC48_113 replaced by BasicMAC48_485

//BasicMAC48_114 replaced by BasicMAC48_485

//BasicMAC48_115 replaced by BasicMAC48_485

//BasicMAC48_116 replaced by BasicMAC48_485

//BasicMAC48_117 replaced by BasicMAC48_485

//BasicMAC48_118 replaced by BasicMAC48_485

//BasicMAC48_119 replaced by BasicMAC48_485

//BasicMAC48_120 replaced by BasicMAC48_485

//BasicMAC48_121 replaced by BasicMAC48_485

//BasicMAC48_122 replaced by BasicMAC48_485

//BasicMAC48_123 replaced by BasicMAC48_485

//BasicMAC48_124 replaced by BasicMAC48_485

//BasicMAC48_125 replaced by BasicMAC48_485

//BasicMAC48_126 replaced by BasicMAC48_485

//BasicMAC48_127 replaced by BasicMAC48_485

//BasicMAC48_128 replaced by BasicMAC48_485

//BasicMAC48_129 replaced by BasicMAC48_485

//BasicMAC48_130 replaced by BasicMAC48_485

//BasicMAC48_131 replaced by BasicMAC48_485

//BasicMAC48_132 replaced by BasicMAC48_485

//BasicMAC48_133 replaced by BasicMAC48_485

//BasicMAC48_134 replaced by BasicMAC48_485

//BasicMAC48_135 replaced by BasicMAC48_485

//BasicMAC48_136 replaced by BasicMAC48_485

//BasicMAC48_137 replaced by BasicMAC48_485

//BasicMAC48_138 replaced by BasicMAC48_485

//BasicMAC48_139 replaced by BasicMAC48_485

//BasicMAC48_140 replaced by BasicMAC48_485

//BasicMAC48_141 replaced by BasicMAC48_485

//BasicMAC48_142 replaced by BasicMAC48_485

//BasicMAC48_143 replaced by BasicMAC48_485

//BasicMAC48_144 replaced by BasicMAC48_485

//BasicMAC48_145 replaced by BasicMAC48_485

//BasicMAC48_146 replaced by BasicMAC48_485

//BasicMAC48_147 replaced by BasicMAC48_485

//BasicMAC48_148 replaced by BasicMAC48_485

//BasicMAC48_149 replaced by BasicMAC48_485

//BasicMAC48_150 replaced by BasicMAC48_485

//BasicMAC48_151 replaced by BasicMAC48_485

//BasicMAC48_152 replaced by BasicMAC48_485

//BasicMAC48_153 replaced by BasicMAC48_485

//BasicMAC48_154 replaced by BasicMAC48_485

//BasicMAC48_155 replaced by BasicMAC48_485

//BasicMAC48_156 replaced by BasicMAC48_485

//BasicMAC48_157 replaced by BasicMAC48_485

//BasicMAC48_158 replaced by BasicMAC48_485

//BasicMAC48_159 replaced by BasicMAC48_485

//BasicMAC48_160 replaced by BasicMAC48_485

//BasicMAC48_161 replaced by BasicMAC48_485

//BasicMAC48_162 replaced by BasicMAC48_485

//BasicMAC48_163 replaced by BasicMAC48_485

//BasicMAC48_164 replaced by BasicMAC48_485

//BasicMAC48_165 replaced by BasicMAC48_485

//BasicMAC48_166 replaced by BasicMAC48_485

//BasicMAC48_167 replaced by BasicMAC48_485

//BasicMAC48_168 replaced by BasicMAC48_485

//BasicMAC48_169 replaced by BasicMAC48_485

//BasicMAC48_170 replaced by BasicMAC48_485

//BasicMAC48_171 replaced by BasicMAC48_485

//BasicMAC48_172 replaced by BasicMAC48_485

//BasicMAC48_173 replaced by BasicMAC48_485

//BasicMAC48_174 replaced by BasicMAC48_485

//BasicMAC48_175 replaced by BasicMAC48_485

//BasicMAC48_176 replaced by BasicMAC48_485

//BasicMAC48_177 replaced by BasicMAC48_485

//BasicMAC48_178 replaced by BasicMAC48_485

//BasicMAC48_179 replaced by BasicMAC48_485

//BasicMAC48_180 replaced by BasicMAC48_485

//BasicMAC48_181 replaced by BasicMAC48_485

//BasicMAC48_182 replaced by BasicMAC48_485

//BasicMAC48_183 replaced by BasicMAC48_485

//BasicMAC48_184 replaced by BasicMAC48_485

//BasicMAC48_185 replaced by BasicMAC48_485

//BasicMAC48_186 replaced by BasicMAC48_485

//BasicMAC48_187 replaced by BasicMAC48_485

//BasicMAC48_188 replaced by BasicMAC48_485

//BasicMAC48_189 replaced by BasicMAC48_485

//BasicMAC48_190 replaced by BasicMAC48_485

//BasicMAC48_191 replaced by BasicMAC48_485

//BasicMAC48_192 replaced by BasicMAC48_485

//BasicMAC48_193 replaced by BasicMAC48_485

//BasicMAC48_194 replaced by BasicMAC48_485

//BasicMAC48_195 replaced by BasicMAC48_485

//BasicMAC48_196 replaced by BasicMAC48_485

//BasicMAC48_197 replaced by BasicMAC48_485

//BasicMAC48_198 replaced by BasicMAC48_485

//BasicMAC48_199 replaced by BasicMAC48_485

//BasicMAC48_200 replaced by BasicMAC48_485

//BasicMAC48_201 replaced by BasicMAC48_485

//BasicMAC48_202 replaced by BasicMAC48_485

//BasicMAC48_203 replaced by BasicMAC48_485

//BasicMAC48_204 replaced by BasicMAC48_485

//BasicMAC48_205 replaced by BasicMAC48_485

//BasicMAC48_206 replaced by BasicMAC48_485

//BasicMAC48_207 replaced by BasicMAC48_485

//BasicMAC48_208 replaced by BasicMAC48_485

//BasicMAC48_209 replaced by BasicMAC48_485

//BasicMAC48_210 replaced by BasicMAC48_485

//BasicMAC48_211 replaced by BasicMAC48_485

//BasicMAC48_212 replaced by BasicMAC48_485

//BasicMAC48_213 replaced by BasicMAC48_485

//BasicMAC48_214 replaced by BasicMAC48_485

//BasicMAC48_215 replaced by BasicMAC48_485

//BasicMAC48_216 replaced by BasicMAC48_485

//BasicMAC48_217 replaced by BasicMAC48_485

//BasicMAC48_218 replaced by BasicMAC48_485

//BasicMAC48_219 replaced by BasicMAC48_485

//BasicMAC48_220 replaced by BasicMAC48_485

//BasicMAC48_221 replaced by BasicMAC48_485

//BasicMAC48_222 replaced by BasicMAC48_485

//BasicMAC48_223 replaced by BasicMAC48_485

//BasicMAC48_224 replaced by BasicMAC48_485

//BasicMAC48_225 replaced by BasicMAC48_485

//BasicMAC48_226 replaced by BasicMAC48_485

//BasicMAC48_227 replaced by BasicMAC48_485

//BasicMAC48_228 replaced by BasicMAC48_485

//BasicMAC48_229 replaced by BasicMAC48_485

//BasicMAC48_230 replaced by BasicMAC48_485

//BasicMAC48_231 replaced by BasicMAC48_485

//BasicMAC48_232 replaced by BasicMAC48_485

//BasicMAC48_233 replaced by BasicMAC48_485

//BasicMAC48_234 replaced by BasicMAC48_485

//BasicMAC48_235 replaced by BasicMAC48_485

//BasicMAC48_236 replaced by BasicMAC48_485

//BasicMAC48_237 replaced by BasicMAC48_485

//BasicMAC48_238 replaced by BasicMAC48_485

//BasicMAC48_239 replaced by BasicMAC48_485

//BasicMAC48_240 replaced by BasicMAC48_485

//BasicMAC48_241 replaced by BasicMAC48_485

//BasicMAC48_242 replaced by BasicMAC48_485

//BasicMAC48_243 replaced by BasicMAC48_485

//BasicMAC48_244 replaced by BasicMAC48_485

//BasicMAC48_245 replaced by BasicMAC48_485

//BasicMAC48_246 replaced by BasicMAC48_485

//BasicMAC48_247 replaced by BasicMAC48_485

//BasicMAC48_248 replaced by BasicMAC48_485

//BasicMAC48_249 replaced by BasicMAC48_485

//BasicMAC48_250 replaced by BasicMAC48_485

//BasicMAC48_251 replaced by BasicMAC48_485

//BasicMAC48_252 replaced by BasicMAC48_485

//BasicMAC48_253 replaced by BasicMAC48_485

//BasicMAC48_254 replaced by BasicMAC48_485

//BasicMAC48_255 replaced by BasicMAC48_485

//BasicMAC48_256 replaced by BasicMAC48_485

//BasicMAC48_257 replaced by BasicMAC48_485

//BasicMAC48_258 replaced by BasicMAC48_485

//BasicMAC48_259 replaced by BasicMAC48_485

//BasicMAC48_260 replaced by BasicMAC48_485

//BasicMAC48_261 replaced by BasicMAC48_485

//BasicMAC48_262 replaced by BasicMAC48_485

//BasicMAC48_263 replaced by BasicMAC48_485

//BasicMAC48_264 replaced by BasicMAC48_485

//BasicMAC48_265 replaced by BasicMAC48_485

//BasicMAC48_266 replaced by BasicMAC48_485

//BasicMAC48_267 replaced by BasicMAC48_485

//BasicMAC48_268 replaced by BasicMAC48_485

//BasicMAC48_269 replaced by BasicMAC48_485

//BasicMAC48_270 replaced by BasicMAC48_485

//BasicMAC48_271 replaced by BasicMAC48_485

//BasicMAC48_272 replaced by BasicMAC48_485

//BasicMAC48_273 replaced by BasicMAC48_485

//BasicMAC48_274 replaced by BasicMAC48_485

//BasicMAC48_275 replaced by BasicMAC48_485

//BasicMAC48_276 replaced by BasicMAC48_485

//BasicMAC48_277 replaced by BasicMAC48_485

//BasicMAC48_278 replaced by BasicMAC48_485

//BasicMAC48_279 replaced by BasicMAC48_485

//BasicMAC48_280 replaced by BasicMAC48_485

//BasicMAC48_281 replaced by BasicMAC48_485

//BasicMAC48_282 replaced by BasicMAC48_485

//BasicMAC48_283 replaced by BasicMAC48_485

//BasicMAC48_284 replaced by BasicMAC48_485

//BasicMAC48_285 replaced by BasicMAC48_485

//BasicMAC48_286 replaced by BasicMAC48_485

//BasicMAC48_287 replaced by BasicMAC48_485

//BasicMAC48_288 replaced by BasicMAC48_485

//BasicMAC48_289 replaced by BasicMAC48_485

//BasicMAC48_290 replaced by BasicMAC48_485

//BasicMAC48_291 replaced by BasicMAC48_485

//BasicMAC48_292 replaced by BasicMAC48_485

//BasicMAC48_293 replaced by BasicMAC48_485

//BasicMAC48_294 replaced by BasicMAC48_485

//BasicMAC48_295 replaced by BasicMAC48_485

//BasicMAC48_296 replaced by BasicMAC48_485

//BasicMAC48_297 replaced by BasicMAC48_485

//BasicMAC48_298 replaced by BasicMAC48_485

//BasicMAC48_299 replaced by BasicMAC48_485

//BasicMAC48_300 replaced by BasicMAC48_485

//BasicMAC48_301 replaced by BasicMAC48_485

//BasicMAC48_302 replaced by BasicMAC48_485

//BasicMAC48_303 replaced by BasicMAC48_485

//BasicMAC48_304 replaced by BasicMAC48_485

//BasicMAC48_305 replaced by BasicMAC48_485

//BasicMAC48_306 replaced by BasicMAC48_485

//BasicMAC48_307 replaced by BasicMAC48_485

//BasicMAC48_308 replaced by BasicMAC48_485

//BasicMAC48_309 replaced by BasicMAC48_485

//BasicMAC48_310 replaced by BasicMAC48_485

//BasicMAC48_311 replaced by BasicMAC48_485

//BasicMAC48_312 replaced by BasicMAC48_485

//BasicMAC48_313 replaced by BasicMAC48_485

//BasicMAC48_314 replaced by BasicMAC48_485

//BasicMAC48_315 replaced by BasicMAC48_485

//BasicMAC48_316 replaced by BasicMAC48_485

//BasicMAC48_317 replaced by BasicMAC48_485

//BasicMAC48_318 replaced by BasicMAC48_485

//BasicMAC48_319 replaced by BasicMAC48_485

//BasicMAC48_320 replaced by BasicMAC48_485

//BasicMAC48_321 replaced by BasicMAC48_485

//BasicMAC48_322 replaced by BasicMAC48_485

//BasicMAC48_323 replaced by BasicMAC48_485

//BasicMAC48_324 replaced by BasicMAC48_485

//BasicMAC48_325 replaced by BasicMAC48_485

//BasicMAC48_326 replaced by BasicMAC48_485

//BasicMAC48_327 replaced by BasicMAC48_485

//BasicMAC48_328 replaced by BasicMAC48_485

//BasicMAC48_329 replaced by BasicMAC48_485

//BasicMAC48_330 replaced by BasicMAC48_485

//BasicMAC48_331 replaced by BasicMAC48_485

//BasicMAC48_332 replaced by BasicMAC48_485

//BasicMAC48_333 replaced by BasicMAC48_485

//BasicMAC48_334 replaced by BasicMAC48_485

//BasicMAC48_335 replaced by BasicMAC48_485

//BasicMAC48_336 replaced by BasicMAC48_485

//BasicMAC48_337 replaced by BasicMAC48_485

//BasicMAC48_338 replaced by BasicMAC48_485

//BasicMAC48_339 replaced by BasicMAC48_485

//BasicMAC48_340 replaced by BasicMAC48_485

//BasicMAC48_341 replaced by BasicMAC48_485

//BasicMAC48_342 replaced by BasicMAC48_485

//BasicMAC48_343 replaced by BasicMAC48_485

//BasicMAC48_344 replaced by BasicMAC48_485

//BasicMAC48_345 replaced by BasicMAC48_485

//BasicMAC48_346 replaced by BasicMAC48_485

//BasicMAC48_347 replaced by BasicMAC48_485

//BasicMAC48_348 replaced by BasicMAC48_485

//BasicMAC48_349 replaced by BasicMAC48_485

//BasicMAC48_350 replaced by BasicMAC48_485

//BasicMAC48_351 replaced by BasicMAC48_485

//BasicMAC48_352 replaced by BasicMAC48_485

//BasicMAC48_353 replaced by BasicMAC48_485

//BasicMAC48_354 replaced by BasicMAC48_485

//BasicMAC48_355 replaced by BasicMAC48_485

//BasicMAC48_356 replaced by BasicMAC48_485

//BasicMAC48_357 replaced by BasicMAC48_485

//BasicMAC48_358 replaced by BasicMAC48_485

//BasicMAC48_359 replaced by BasicMAC48_485

//BasicMAC48_360 replaced by BasicMAC48_485

//BasicMAC48_361 replaced by BasicMAC48_485

//BasicMAC48_362 replaced by BasicMAC48_485

//BasicMAC48_363 replaced by BasicMAC48_485

//BasicMAC48_364 replaced by BasicMAC48_485

//BasicMAC48_365 replaced by BasicMAC48_485

//BasicMAC48_366 replaced by BasicMAC48_485

//BasicMAC48_367 replaced by BasicMAC48_485

//BasicMAC48_368 replaced by BasicMAC48_485

//BasicMAC48_369 replaced by BasicMAC48_485

//BasicMAC48_370 replaced by BasicMAC48_485

//BasicMAC48_371 replaced by BasicMAC48_485

//BasicMAC48_372 replaced by BasicMAC48_485

//BasicMAC48_373 replaced by BasicMAC48_485

//BasicMAC48_374 replaced by BasicMAC48_485

//BasicMAC48_375 replaced by BasicMAC48_485

//BasicMAC48_376 replaced by BasicMAC48_485

//BasicMAC48_377 replaced by BasicMAC48_485

//BasicMAC48_378 replaced by BasicMAC48_485

//BasicMAC48_379 replaced by BasicMAC48_485

//BasicMAC48_380 replaced by BasicMAC48_485

//BasicMAC48_381 replaced by BasicMAC48_485

//BasicMAC48_382 replaced by BasicMAC48_485

//BasicMAC48_383 replaced by BasicMAC48_485

//BasicMAC48_384 replaced by BasicMAC48_485

//BasicMAC48_385 replaced by BasicMAC48_485

//BasicMAC48_386 replaced by BasicMAC48_485

//BasicMAC48_387 replaced by BasicMAC48_485

//BasicMAC48_388 replaced by BasicMAC48_485

//BasicMAC48_389 replaced by BasicMAC48_485

//BasicMAC48_390 replaced by BasicMAC48_485

//BasicMAC48_391 replaced by BasicMAC48_485

//BasicMAC48_392 replaced by BasicMAC48_485

//BasicMAC48_393 replaced by BasicMAC48_485

//BasicMAC48_394 replaced by BasicMAC48_485

//BasicMAC48_395 replaced by BasicMAC48_485

//BasicMAC48_396 replaced by BasicMAC48_485

//BasicMAC48_397 replaced by BasicMAC48_485

//BasicMAC48_398 replaced by BasicMAC48_485

//BasicMAC48_399 replaced by BasicMAC48_485

//BasicMAC48_400 replaced by BasicMAC48_485

//BasicMAC48_401 replaced by BasicMAC48_485

//BasicMAC48_402 replaced by BasicMAC48_485

//BasicMAC48_403 replaced by BasicMAC48_485

//BasicMAC48_404 replaced by BasicMAC48_485

//BasicMAC48_405 replaced by BasicMAC48_485

//BasicMAC48_406 replaced by BasicMAC48_485

//BasicMAC48_407 replaced by BasicMAC48_485

//BasicMAC48_408 replaced by BasicMAC48_485

//BasicMAC48_409 replaced by BasicMAC48_485

//BasicMAC48_410 replaced by BasicMAC48_485

//BasicMAC48_411 replaced by BasicMAC48_485

//BasicMAC48_412 replaced by BasicMAC48_485

//BasicMAC48_413 replaced by BasicMAC48_485

//BasicMAC48_414 replaced by BasicMAC48_485

//BasicMAC48_415 replaced by BasicMAC48_485

//BasicMAC48_416 replaced by BasicMAC48_485

//BasicMAC48_417 replaced by BasicMAC48_485

//BasicMAC48_418 replaced by BasicMAC48_485

//BasicMAC48_419 replaced by BasicMAC48_485

//BasicMAC48_420 replaced by BasicMAC48_485

//BasicMAC48_421 replaced by BasicMAC48_485

//BasicMAC48_422 replaced by BasicMAC48_485

//BasicMAC48_423 replaced by BasicMAC48_485

//BasicMAC48_424 replaced by BasicMAC48_485

//BasicMAC48_425 replaced by BasicMAC48_485

//BasicMAC48_426 replaced by BasicMAC48_485

//BasicMAC48_427 replaced by BasicMAC48_485

//BasicMAC48_428 replaced by BasicMAC48_485

//BasicMAC48_429 replaced by BasicMAC48_485

//BasicMAC48_430 replaced by BasicMAC48_485

//BasicMAC48_431 replaced by BasicMAC48_485

//BasicMAC48_432 replaced by BasicMAC48_485

//BasicMAC48_433 replaced by BasicMAC48_485

//BasicMAC48_434 replaced by BasicMAC48_485

//BasicMAC48_435 replaced by BasicMAC48_485

//BasicMAC48_436 replaced by BasicMAC48_485

//BasicMAC48_437 replaced by BasicMAC48_485

//BasicMAC48_438 replaced by BasicMAC48_485

//BasicMAC48_439 replaced by BasicMAC48_485

//BasicMAC48_440 replaced by BasicMAC48_485

//BasicMAC48_441 replaced by BasicMAC48_485

//BasicMAC48_442 replaced by BasicMAC48_485

//BasicMAC48_443 replaced by BasicMAC48_485

//BasicMAC48_444 replaced by BasicMAC48_485

//BasicMAC48_445 replaced by BasicMAC48_485

//BasicMAC48_446 replaced by BasicMAC48_485

//BasicMAC48_447 replaced by BasicMAC48_485

//BasicMAC48_448 replaced by BasicMAC48_485

//BasicMAC48_449 replaced by BasicMAC48_485

//BasicMAC48_450 replaced by BasicMAC48_485

//BasicMAC48_451 replaced by BasicMAC48_485

//BasicMAC48_452 replaced by BasicMAC48_485

//BasicMAC48_453 replaced by BasicMAC48_485

//BasicMAC48_454 replaced by BasicMAC48_485

//BasicMAC48_455 replaced by BasicMAC48_485

//BasicMAC48_456 replaced by BasicMAC48_485

//BasicMAC48_457 replaced by BasicMAC48_485

//BasicMAC48_458 replaced by BasicMAC48_485

//BasicMAC48_459 replaced by BasicMAC48_485

//BasicMAC48_460 replaced by BasicMAC48_485

//BasicMAC48_461 replaced by BasicMAC48_485

//BasicMAC48_462 replaced by BasicMAC48_485

//BasicMAC48_463 replaced by BasicMAC48_485

//BasicMAC48_464 replaced by BasicMAC48_485

//BasicMAC48_465 replaced by BasicMAC48_485

//BasicMAC48_466 replaced by BasicMAC48_485

//BasicMAC48_467 replaced by BasicMAC48_485

//BasicMAC48_468 replaced by BasicMAC48_485

//BasicMAC48_469 replaced by BasicMAC48_485

//BasicMAC48_470 replaced by BasicMAC48_485

//BasicMAC48_471 replaced by BasicMAC48_485

//BasicMAC48_472 replaced by BasicMAC48_485

//BasicMAC48_473 replaced by BasicMAC48_485

//BasicMAC48_474 replaced by BasicMAC48_485

//BasicMAC48_475 replaced by BasicMAC48_485

//BasicMAC48_476 replaced by BasicMAC48_485

//BasicMAC48_477 replaced by BasicMAC48_485

//BasicMAC48_478 replaced by BasicMAC48_485

//BasicMAC48_479 replaced by BasicMAC48_485

//BasicMAC48_480 replaced by BasicMAC48_485

//BasicMAC48_481 replaced by BasicMAC48_485

//BasicMAC48_482 replaced by BasicMAC48_485

//BasicMAC48_483 replaced by BasicMAC48_485

//BasicMAC48_484 replaced by BasicMAC48_485

module BasicMAC48_485 (
  input      [51:0]   io_a,
  input      [50:0]   io_b,
  input      [50:0]   io_c,
  input               io_ce,
  output reg [102:0]  io_p,
  input               clk,
  input               resetn
);

  wire       [25:0]   MACs_0_0_io_a;
  wire       [16:0]   MACs_0_0_io_b;
  reg        [16:0]   MACs_1_0_io_c;
  wire       [29:0]   MACs_0_0_io_acout;
  wire       [42:0]   MACs_0_0_io_p;
  wire       [47:0]   MACs_0_0_io_pcout;
  wire       [29:0]   MACs_0_1_io_acout;
  wire       [42:0]   MACs_0_1_io_p;
  wire       [47:0]   MACs_0_1_io_pcout;
  wire       [29:0]   MACs_0_2_io_acout;
  wire       [42:0]   MACs_0_2_io_p;
  wire       [47:0]   MACs_0_2_io_pcout;
  wire       [29:0]   MACs_1_0_io_acout;
  wire       [42:0]   MACs_1_0_io_p;
  wire       [47:0]   MACs_1_0_io_pcout;
  wire       [29:0]   MACs_1_1_io_acout;
  wire       [42:0]   MACs_1_1_io_p;
  wire       [47:0]   MACs_1_1_io_pcout;
  wire       [29:0]   MACs_1_2_io_acout;
  wire       [42:0]   MACs_1_2_io_p;
  wire       [47:0]   MACs_1_2_io_pcout;
  reg        [16:0]   _zz_io_b;
  reg        [16:0]   _zz_io_b_1;
  reg        [16:0]   _zz_io_b_2;
  reg        [16:0]   _zz_io_c;
  reg        [16:0]   _zz_io_c_1;
  reg        [16:0]   _zz_io_c_2;
  reg        [16:0]   _zz_io_c_3;
  reg        [16:0]   _zz_io_c_4;
  reg        [16:0]   _zz_io_c_5;
  reg                 _zz_io_ce;
  reg                 _zz_io_ce_1;
  reg                 _zz_io_ce_2;
  reg        [25:0]   _zz_io_a;
  reg        [25:0]   _zz_io_a_1;
  reg        [25:0]   _zz_io_a_2;
  reg        [25:0]   _zz_io_a_3;
  reg        [16:0]   _zz_io_b_3;
  reg        [16:0]   _zz_io_b_4;
  reg        [16:0]   _zz_io_b_5;
  reg        [16:0]   _zz_io_b_6;
  reg        [16:0]   _zz_io_b_7;
  reg        [16:0]   _zz_io_b_8;
  reg        [16:0]   _zz_io_b_9;
  reg        [16:0]   _zz_io_b_10;
  reg        [16:0]   _zz_io_b_11;
  reg        [16:0]   _zz_io_b_12;
  reg        [16:0]   _zz_io_b_13;
  reg        [16:0]   _zz_io_b_14;
  reg        [7:0]    _zz_io_c_6;
  reg        [16:0]   _zz_io_c_7;
  reg        [16:0]   _zz_io_c_8;
  reg        [16:0]   _zz_io_c_9;
  reg        [16:0]   _zz_io_p;
  reg        [16:0]   _zz_io_p_1;
  reg        [16:0]   _zz_io_p_2;
  reg        [16:0]   _zz_io_p_3;
  reg        [16:0]   _zz_io_p_4;
  reg        [8:0]    _zz_io_p_5;
  reg        [8:0]    _zz_io_p_6;
  reg        [8:0]    _zz_io_p_7;
  reg        [8:0]    _zz_io_p_8;
  reg        [16:0]   _zz_io_p_9;
  reg        [11:0]   _zz_io_p_10;
  reg        [6:0]    _zz_io_p_11;

  MAC_2910 MACs_0_0 (
    .io_a     (MACs_0_0_io_a[25:0]    ), //i
    .io_acin  (30'h0                  ), //i
    .io_acout (MACs_0_0_io_acout[29:0]), //o
    .io_b     (MACs_0_0_io_b[16:0]    ), //i
    .io_c     (_zz_io_c[16:0]         ), //i
    .io_ce    (_zz_io_ce              ), //i
    .io_pcin  (48'h0                  ), //i
    .io_p     (MACs_0_0_io_p[42:0]    ), //o
    .io_pcout (MACs_0_0_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_2911 MACs_0_1 (
    .io_a     (26'h0                  ), //i
    .io_acin  (MACs_0_0_io_acout[29:0]), //i
    .io_acout (MACs_0_1_io_acout[29:0]), //o
    .io_b     (_zz_io_b[16:0]         ), //i
    .io_c     (_zz_io_c_2[16:0]       ), //i
    .io_ce    (_zz_io_ce_1            ), //i
    .io_pcin  (MACs_0_0_io_pcout[47:0]), //i
    .io_p     (MACs_0_1_io_p[42:0]    ), //o
    .io_pcout (MACs_0_1_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_2911 MACs_0_2 (
    .io_a     (26'h0                  ), //i
    .io_acin  (MACs_0_1_io_acout[29:0]), //i
    .io_acout (MACs_0_2_io_acout[29:0]), //o
    .io_b     (_zz_io_b_2[16:0]       ), //i
    .io_c     (_zz_io_c_5[16:0]       ), //i
    .io_ce    (_zz_io_ce_2            ), //i
    .io_pcin  (MACs_0_1_io_pcout[47:0]), //i
    .io_p     (MACs_0_2_io_p[42:0]    ), //o
    .io_pcout (MACs_0_2_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_2910 MACs_1_0 (
    .io_a     (_zz_io_a_3[25:0]       ), //i
    .io_acin  (30'h0                  ), //i
    .io_acout (MACs_1_0_io_acout[29:0]), //o
    .io_b     (_zz_io_b_12[16:0]      ), //i
    .io_c     (MACs_1_0_io_c[16:0]    ), //i
    .io_ce    (1'b1                   ), //i
    .io_pcin  (48'h0                  ), //i
    .io_p     (MACs_1_0_io_p[42:0]    ), //o
    .io_pcout (MACs_1_0_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_2911 MACs_1_1 (
    .io_a     (26'h0                  ), //i
    .io_acin  (MACs_1_0_io_acout[29:0]), //i
    .io_acout (MACs_1_1_io_acout[29:0]), //o
    .io_b     (_zz_io_b_13[16:0]      ), //i
    .io_c     (_zz_io_c_7[16:0]       ), //i
    .io_ce    (1'b1                   ), //i
    .io_pcin  (MACs_1_0_io_pcout[47:0]), //i
    .io_p     (MACs_1_1_io_p[42:0]    ), //o
    .io_pcout (MACs_1_1_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  MAC_2911 MACs_1_2 (
    .io_a     (26'h0                  ), //i
    .io_acin  (MACs_1_1_io_acout[29:0]), //i
    .io_acout (MACs_1_2_io_acout[29:0]), //o
    .io_b     (_zz_io_b_14[16:0]      ), //i
    .io_c     (_zz_io_c_9[16:0]       ), //i
    .io_ce    (1'b1                   ), //i
    .io_pcin  (MACs_1_1_io_pcout[47:0]), //i
    .io_p     (MACs_1_2_io_p[42:0]    ), //o
    .io_pcout (MACs_1_2_io_pcout[47:0]), //o
    .clk      (clk                    )  //i
  );
  assign MACs_0_0_io_a = io_a[25:0];
  assign MACs_0_0_io_b = io_b[16 : 0];
  always @(*) begin
    MACs_1_0_io_c[7 : 0] = _zz_io_c_6;
    MACs_1_0_io_c[16 : 8] = MACs_0_2_io_p[8 : 0];
  end

  always @(*) begin
    io_p[16 : 0] = _zz_io_p_4;
    io_p[25 : 17] = _zz_io_p_8;
    io_p[42 : 26] = _zz_io_p_9;
    io_p[47 : 43] = MACs_1_1_io_p[4 : 0];
    io_p[59 : 48] = _zz_io_p_10;
    io_p[95 : 60] = MACs_1_2_io_p[35 : 0];
    io_p[102 : 96] = _zz_io_p_11;
  end

  always @(posedge clk) begin
    _zz_io_b <= io_b[33 : 17];
    _zz_io_b_1 <= io_b[50 : 34];
    _zz_io_b_2 <= _zz_io_b_1;
    _zz_io_c <= io_c[16 : 0];
    _zz_io_c_1 <= io_c[33 : 17];
    _zz_io_c_2 <= _zz_io_c_1;
    _zz_io_c_3 <= io_c[50 : 34];
    _zz_io_c_4 <= _zz_io_c_3;
    _zz_io_c_5 <= _zz_io_c_4;
    _zz_io_ce <= io_ce;
    _zz_io_ce_1 <= _zz_io_ce;
    _zz_io_ce_2 <= _zz_io_ce_1;
    _zz_io_a <= (io_a >>> 26);
    _zz_io_a_1 <= _zz_io_a;
    _zz_io_a_2 <= _zz_io_a_1;
    _zz_io_a_3 <= _zz_io_a_2;
    _zz_io_b_3 <= MACs_0_0_io_b;
    _zz_io_b_4 <= _zz_io_b;
    _zz_io_b_5 <= _zz_io_b_2;
    _zz_io_b_6 <= _zz_io_b_3;
    _zz_io_b_7 <= _zz_io_b_4;
    _zz_io_b_8 <= _zz_io_b_5;
    _zz_io_b_9 <= _zz_io_b_6;
    _zz_io_b_10 <= _zz_io_b_7;
    _zz_io_b_11 <= _zz_io_b_8;
    _zz_io_b_12 <= _zz_io_b_9;
    _zz_io_b_13 <= _zz_io_b_10;
    _zz_io_b_14 <= _zz_io_b_11;
    _zz_io_c_6 <= MACs_0_1_io_p[16 : 9];
    _zz_io_c_7 <= MACs_0_2_io_p[25 : 9];
    _zz_io_c_8 <= MACs_0_2_io_p[42 : 26];
    _zz_io_c_9 <= _zz_io_c_8;
    _zz_io_p <= MACs_0_0_io_p[16 : 0];
    _zz_io_p_1 <= _zz_io_p;
    _zz_io_p_2 <= _zz_io_p_1;
    _zz_io_p_3 <= _zz_io_p_2;
    _zz_io_p_4 <= _zz_io_p_3;
    _zz_io_p_5 <= MACs_0_1_io_p[8 : 0];
    _zz_io_p_6 <= _zz_io_p_5;
    _zz_io_p_7 <= _zz_io_p_6;
    _zz_io_p_8 <= _zz_io_p_7;
    _zz_io_p_9 <= MACs_1_0_io_p[16 : 0];
    _zz_io_p_10 <= MACs_1_1_io_p[16 : 5];
    _zz_io_p_11 <= MACs_1_2_io_p[42 : 36];
  end


endmodule

//MAC_5 replaced by MAC_2911

//MAC_4 replaced by MAC_2911

//MAC_3 replaced by MAC_2910

//MAC_2 replaced by MAC_2911

//MAC_1 replaced by MAC_2911

//MAC replaced by MAC_2910

//MAC_11 replaced by MAC_2911

//MAC_10 replaced by MAC_2911

//MAC_9 replaced by MAC_2910

//MAC_8 replaced by MAC_2911

//MAC_7 replaced by MAC_2911

//MAC_6 replaced by MAC_2910

//MAC_17 replaced by MAC_2911

//MAC_16 replaced by MAC_2911

//MAC_15 replaced by MAC_2910

//MAC_14 replaced by MAC_2911

//MAC_13 replaced by MAC_2911

//MAC_12 replaced by MAC_2910

//MAC_23 replaced by MAC_2911

//MAC_22 replaced by MAC_2911

//MAC_21 replaced by MAC_2910

//MAC_20 replaced by MAC_2911

//MAC_19 replaced by MAC_2911

//MAC_18 replaced by MAC_2910

//MAC_29 replaced by MAC_2911

//MAC_28 replaced by MAC_2911

//MAC_27 replaced by MAC_2910

//MAC_26 replaced by MAC_2911

//MAC_25 replaced by MAC_2911

//MAC_24 replaced by MAC_2910

//MAC_35 replaced by MAC_2911

//MAC_34 replaced by MAC_2911

//MAC_33 replaced by MAC_2910

//MAC_32 replaced by MAC_2911

//MAC_31 replaced by MAC_2911

//MAC_30 replaced by MAC_2910

//MAC_41 replaced by MAC_2911

//MAC_40 replaced by MAC_2911

//MAC_39 replaced by MAC_2910

//MAC_38 replaced by MAC_2911

//MAC_37 replaced by MAC_2911

//MAC_36 replaced by MAC_2910

//MAC_47 replaced by MAC_2911

//MAC_46 replaced by MAC_2911

//MAC_45 replaced by MAC_2910

//MAC_44 replaced by MAC_2911

//MAC_43 replaced by MAC_2911

//MAC_42 replaced by MAC_2910

//MAC_53 replaced by MAC_2911

//MAC_52 replaced by MAC_2911

//MAC_51 replaced by MAC_2910

//MAC_50 replaced by MAC_2911

//MAC_49 replaced by MAC_2911

//MAC_48 replaced by MAC_2910

//MAC_59 replaced by MAC_2911

//MAC_58 replaced by MAC_2911

//MAC_57 replaced by MAC_2910

//MAC_56 replaced by MAC_2911

//MAC_55 replaced by MAC_2911

//MAC_54 replaced by MAC_2910

//MAC_65 replaced by MAC_2911

//MAC_64 replaced by MAC_2911

//MAC_63 replaced by MAC_2910

//MAC_62 replaced by MAC_2911

//MAC_61 replaced by MAC_2911

//MAC_60 replaced by MAC_2910

//MAC_71 replaced by MAC_2911

//MAC_70 replaced by MAC_2911

//MAC_69 replaced by MAC_2910

//MAC_68 replaced by MAC_2911

//MAC_67 replaced by MAC_2911

//MAC_66 replaced by MAC_2910

//MAC_77 replaced by MAC_2911

//MAC_76 replaced by MAC_2911

//MAC_75 replaced by MAC_2910

//MAC_74 replaced by MAC_2911

//MAC_73 replaced by MAC_2911

//MAC_72 replaced by MAC_2910

//MAC_83 replaced by MAC_2911

//MAC_82 replaced by MAC_2911

//MAC_81 replaced by MAC_2910

//MAC_80 replaced by MAC_2911

//MAC_79 replaced by MAC_2911

//MAC_78 replaced by MAC_2910

//MAC_89 replaced by MAC_2911

//MAC_88 replaced by MAC_2911

//MAC_87 replaced by MAC_2910

//MAC_86 replaced by MAC_2911

//MAC_85 replaced by MAC_2911

//MAC_84 replaced by MAC_2910

//MAC_95 replaced by MAC_2911

//MAC_94 replaced by MAC_2911

//MAC_93 replaced by MAC_2910

//MAC_92 replaced by MAC_2911

//MAC_91 replaced by MAC_2911

//MAC_90 replaced by MAC_2910

//MAC_101 replaced by MAC_2911

//MAC_100 replaced by MAC_2911

//MAC_99 replaced by MAC_2910

//MAC_98 replaced by MAC_2911

//MAC_97 replaced by MAC_2911

//MAC_96 replaced by MAC_2910

//MAC_107 replaced by MAC_2911

//MAC_106 replaced by MAC_2911

//MAC_105 replaced by MAC_2910

//MAC_104 replaced by MAC_2911

//MAC_103 replaced by MAC_2911

//MAC_102 replaced by MAC_2910

//MAC_113 replaced by MAC_2911

//MAC_112 replaced by MAC_2911

//MAC_111 replaced by MAC_2910

//MAC_110 replaced by MAC_2911

//MAC_109 replaced by MAC_2911

//MAC_108 replaced by MAC_2910

//MAC_119 replaced by MAC_2911

//MAC_118 replaced by MAC_2911

//MAC_117 replaced by MAC_2910

//MAC_116 replaced by MAC_2911

//MAC_115 replaced by MAC_2911

//MAC_114 replaced by MAC_2910

//MAC_125 replaced by MAC_2911

//MAC_124 replaced by MAC_2911

//MAC_123 replaced by MAC_2910

//MAC_122 replaced by MAC_2911

//MAC_121 replaced by MAC_2911

//MAC_120 replaced by MAC_2910

//MAC_131 replaced by MAC_2911

//MAC_130 replaced by MAC_2911

//MAC_129 replaced by MAC_2910

//MAC_128 replaced by MAC_2911

//MAC_127 replaced by MAC_2911

//MAC_126 replaced by MAC_2910

//MAC_137 replaced by MAC_2911

//MAC_136 replaced by MAC_2911

//MAC_135 replaced by MAC_2910

//MAC_134 replaced by MAC_2911

//MAC_133 replaced by MAC_2911

//MAC_132 replaced by MAC_2910

//MAC_143 replaced by MAC_2911

//MAC_142 replaced by MAC_2911

//MAC_141 replaced by MAC_2910

//MAC_140 replaced by MAC_2911

//MAC_139 replaced by MAC_2911

//MAC_138 replaced by MAC_2910

//MAC_149 replaced by MAC_2911

//MAC_148 replaced by MAC_2911

//MAC_147 replaced by MAC_2910

//MAC_146 replaced by MAC_2911

//MAC_145 replaced by MAC_2911

//MAC_144 replaced by MAC_2910

//MAC_155 replaced by MAC_2911

//MAC_154 replaced by MAC_2911

//MAC_153 replaced by MAC_2910

//MAC_152 replaced by MAC_2911

//MAC_151 replaced by MAC_2911

//MAC_150 replaced by MAC_2910

//MAC_161 replaced by MAC_2911

//MAC_160 replaced by MAC_2911

//MAC_159 replaced by MAC_2910

//MAC_158 replaced by MAC_2911

//MAC_157 replaced by MAC_2911

//MAC_156 replaced by MAC_2910

//MAC_167 replaced by MAC_2911

//MAC_166 replaced by MAC_2911

//MAC_165 replaced by MAC_2910

//MAC_164 replaced by MAC_2911

//MAC_163 replaced by MAC_2911

//MAC_162 replaced by MAC_2910

//MAC_173 replaced by MAC_2911

//MAC_172 replaced by MAC_2911

//MAC_171 replaced by MAC_2910

//MAC_170 replaced by MAC_2911

//MAC_169 replaced by MAC_2911

//MAC_168 replaced by MAC_2910

//MAC_179 replaced by MAC_2911

//MAC_178 replaced by MAC_2911

//MAC_177 replaced by MAC_2910

//MAC_176 replaced by MAC_2911

//MAC_175 replaced by MAC_2911

//MAC_174 replaced by MAC_2910

//MAC_185 replaced by MAC_2911

//MAC_184 replaced by MAC_2911

//MAC_183 replaced by MAC_2910

//MAC_182 replaced by MAC_2911

//MAC_181 replaced by MAC_2911

//MAC_180 replaced by MAC_2910

//MAC_191 replaced by MAC_2911

//MAC_190 replaced by MAC_2911

//MAC_189 replaced by MAC_2910

//MAC_188 replaced by MAC_2911

//MAC_187 replaced by MAC_2911

//MAC_186 replaced by MAC_2910

//MAC_197 replaced by MAC_2911

//MAC_196 replaced by MAC_2911

//MAC_195 replaced by MAC_2910

//MAC_194 replaced by MAC_2911

//MAC_193 replaced by MAC_2911

//MAC_192 replaced by MAC_2910

//MAC_203 replaced by MAC_2911

//MAC_202 replaced by MAC_2911

//MAC_201 replaced by MAC_2910

//MAC_200 replaced by MAC_2911

//MAC_199 replaced by MAC_2911

//MAC_198 replaced by MAC_2910

//MAC_209 replaced by MAC_2911

//MAC_208 replaced by MAC_2911

//MAC_207 replaced by MAC_2910

//MAC_206 replaced by MAC_2911

//MAC_205 replaced by MAC_2911

//MAC_204 replaced by MAC_2910

//MAC_215 replaced by MAC_2911

//MAC_214 replaced by MAC_2911

//MAC_213 replaced by MAC_2910

//MAC_212 replaced by MAC_2911

//MAC_211 replaced by MAC_2911

//MAC_210 replaced by MAC_2910

//MAC_221 replaced by MAC_2911

//MAC_220 replaced by MAC_2911

//MAC_219 replaced by MAC_2910

//MAC_218 replaced by MAC_2911

//MAC_217 replaced by MAC_2911

//MAC_216 replaced by MAC_2910

//MAC_227 replaced by MAC_2911

//MAC_226 replaced by MAC_2911

//MAC_225 replaced by MAC_2910

//MAC_224 replaced by MAC_2911

//MAC_223 replaced by MAC_2911

//MAC_222 replaced by MAC_2910

//MAC_233 replaced by MAC_2911

//MAC_232 replaced by MAC_2911

//MAC_231 replaced by MAC_2910

//MAC_230 replaced by MAC_2911

//MAC_229 replaced by MAC_2911

//MAC_228 replaced by MAC_2910

//MAC_239 replaced by MAC_2911

//MAC_238 replaced by MAC_2911

//MAC_237 replaced by MAC_2910

//MAC_236 replaced by MAC_2911

//MAC_235 replaced by MAC_2911

//MAC_234 replaced by MAC_2910

//MAC_245 replaced by MAC_2911

//MAC_244 replaced by MAC_2911

//MAC_243 replaced by MAC_2910

//MAC_242 replaced by MAC_2911

//MAC_241 replaced by MAC_2911

//MAC_240 replaced by MAC_2910

//MAC_251 replaced by MAC_2911

//MAC_250 replaced by MAC_2911

//MAC_249 replaced by MAC_2910

//MAC_248 replaced by MAC_2911

//MAC_247 replaced by MAC_2911

//MAC_246 replaced by MAC_2910

//MAC_257 replaced by MAC_2911

//MAC_256 replaced by MAC_2911

//MAC_255 replaced by MAC_2910

//MAC_254 replaced by MAC_2911

//MAC_253 replaced by MAC_2911

//MAC_252 replaced by MAC_2910

//MAC_263 replaced by MAC_2911

//MAC_262 replaced by MAC_2911

//MAC_261 replaced by MAC_2910

//MAC_260 replaced by MAC_2911

//MAC_259 replaced by MAC_2911

//MAC_258 replaced by MAC_2910

//MAC_269 replaced by MAC_2911

//MAC_268 replaced by MAC_2911

//MAC_267 replaced by MAC_2910

//MAC_266 replaced by MAC_2911

//MAC_265 replaced by MAC_2911

//MAC_264 replaced by MAC_2910

//MAC_275 replaced by MAC_2911

//MAC_274 replaced by MAC_2911

//MAC_273 replaced by MAC_2910

//MAC_272 replaced by MAC_2911

//MAC_271 replaced by MAC_2911

//MAC_270 replaced by MAC_2910

//MAC_281 replaced by MAC_2911

//MAC_280 replaced by MAC_2911

//MAC_279 replaced by MAC_2910

//MAC_278 replaced by MAC_2911

//MAC_277 replaced by MAC_2911

//MAC_276 replaced by MAC_2910

//MAC_287 replaced by MAC_2911

//MAC_286 replaced by MAC_2911

//MAC_285 replaced by MAC_2910

//MAC_284 replaced by MAC_2911

//MAC_283 replaced by MAC_2911

//MAC_282 replaced by MAC_2910

//MAC_293 replaced by MAC_2911

//MAC_292 replaced by MAC_2911

//MAC_291 replaced by MAC_2910

//MAC_290 replaced by MAC_2911

//MAC_289 replaced by MAC_2911

//MAC_288 replaced by MAC_2910

//MAC_299 replaced by MAC_2911

//MAC_298 replaced by MAC_2911

//MAC_297 replaced by MAC_2910

//MAC_296 replaced by MAC_2911

//MAC_295 replaced by MAC_2911

//MAC_294 replaced by MAC_2910

//MAC_305 replaced by MAC_2911

//MAC_304 replaced by MAC_2911

//MAC_303 replaced by MAC_2910

//MAC_302 replaced by MAC_2911

//MAC_301 replaced by MAC_2911

//MAC_300 replaced by MAC_2910

//MAC_311 replaced by MAC_2911

//MAC_310 replaced by MAC_2911

//MAC_309 replaced by MAC_2910

//MAC_308 replaced by MAC_2911

//MAC_307 replaced by MAC_2911

//MAC_306 replaced by MAC_2910

//MAC_317 replaced by MAC_2911

//MAC_316 replaced by MAC_2911

//MAC_315 replaced by MAC_2910

//MAC_314 replaced by MAC_2911

//MAC_313 replaced by MAC_2911

//MAC_312 replaced by MAC_2910

//MAC_323 replaced by MAC_2911

//MAC_322 replaced by MAC_2911

//MAC_321 replaced by MAC_2910

//MAC_320 replaced by MAC_2911

//MAC_319 replaced by MAC_2911

//MAC_318 replaced by MAC_2910

//MAC_329 replaced by MAC_2911

//MAC_328 replaced by MAC_2911

//MAC_327 replaced by MAC_2910

//MAC_326 replaced by MAC_2911

//MAC_325 replaced by MAC_2911

//MAC_324 replaced by MAC_2910

//MAC_335 replaced by MAC_2911

//MAC_334 replaced by MAC_2911

//MAC_333 replaced by MAC_2910

//MAC_332 replaced by MAC_2911

//MAC_331 replaced by MAC_2911

//MAC_330 replaced by MAC_2910

//MAC_341 replaced by MAC_2911

//MAC_340 replaced by MAC_2911

//MAC_339 replaced by MAC_2910

//MAC_338 replaced by MAC_2911

//MAC_337 replaced by MAC_2911

//MAC_336 replaced by MAC_2910

//MAC_347 replaced by MAC_2911

//MAC_346 replaced by MAC_2911

//MAC_345 replaced by MAC_2910

//MAC_344 replaced by MAC_2911

//MAC_343 replaced by MAC_2911

//MAC_342 replaced by MAC_2910

//MAC_353 replaced by MAC_2911

//MAC_352 replaced by MAC_2911

//MAC_351 replaced by MAC_2910

//MAC_350 replaced by MAC_2911

//MAC_349 replaced by MAC_2911

//MAC_348 replaced by MAC_2910

//MAC_359 replaced by MAC_2911

//MAC_358 replaced by MAC_2911

//MAC_357 replaced by MAC_2910

//MAC_356 replaced by MAC_2911

//MAC_355 replaced by MAC_2911

//MAC_354 replaced by MAC_2910

//MAC_365 replaced by MAC_2911

//MAC_364 replaced by MAC_2911

//MAC_363 replaced by MAC_2910

//MAC_362 replaced by MAC_2911

//MAC_361 replaced by MAC_2911

//MAC_360 replaced by MAC_2910

//MAC_371 replaced by MAC_2911

//MAC_370 replaced by MAC_2911

//MAC_369 replaced by MAC_2910

//MAC_368 replaced by MAC_2911

//MAC_367 replaced by MAC_2911

//MAC_366 replaced by MAC_2910

//MAC_377 replaced by MAC_2911

//MAC_376 replaced by MAC_2911

//MAC_375 replaced by MAC_2910

//MAC_374 replaced by MAC_2911

//MAC_373 replaced by MAC_2911

//MAC_372 replaced by MAC_2910

//MAC_383 replaced by MAC_2911

//MAC_382 replaced by MAC_2911

//MAC_381 replaced by MAC_2910

//MAC_380 replaced by MAC_2911

//MAC_379 replaced by MAC_2911

//MAC_378 replaced by MAC_2910

//MAC_389 replaced by MAC_2911

//MAC_388 replaced by MAC_2911

//MAC_387 replaced by MAC_2910

//MAC_386 replaced by MAC_2911

//MAC_385 replaced by MAC_2911

//MAC_384 replaced by MAC_2910

//MAC_395 replaced by MAC_2911

//MAC_394 replaced by MAC_2911

//MAC_393 replaced by MAC_2910

//MAC_392 replaced by MAC_2911

//MAC_391 replaced by MAC_2911

//MAC_390 replaced by MAC_2910

//MAC_401 replaced by MAC_2911

//MAC_400 replaced by MAC_2911

//MAC_399 replaced by MAC_2910

//MAC_398 replaced by MAC_2911

//MAC_397 replaced by MAC_2911

//MAC_396 replaced by MAC_2910

//MAC_407 replaced by MAC_2911

//MAC_406 replaced by MAC_2911

//MAC_405 replaced by MAC_2910

//MAC_404 replaced by MAC_2911

//MAC_403 replaced by MAC_2911

//MAC_402 replaced by MAC_2910

//MAC_413 replaced by MAC_2911

//MAC_412 replaced by MAC_2911

//MAC_411 replaced by MAC_2910

//MAC_410 replaced by MAC_2911

//MAC_409 replaced by MAC_2911

//MAC_408 replaced by MAC_2910

//MAC_419 replaced by MAC_2911

//MAC_418 replaced by MAC_2911

//MAC_417 replaced by MAC_2910

//MAC_416 replaced by MAC_2911

//MAC_415 replaced by MAC_2911

//MAC_414 replaced by MAC_2910

//MAC_425 replaced by MAC_2911

//MAC_424 replaced by MAC_2911

//MAC_423 replaced by MAC_2910

//MAC_422 replaced by MAC_2911

//MAC_421 replaced by MAC_2911

//MAC_420 replaced by MAC_2910

//MAC_431 replaced by MAC_2911

//MAC_430 replaced by MAC_2911

//MAC_429 replaced by MAC_2910

//MAC_428 replaced by MAC_2911

//MAC_427 replaced by MAC_2911

//MAC_426 replaced by MAC_2910

//MAC_437 replaced by MAC_2911

//MAC_436 replaced by MAC_2911

//MAC_435 replaced by MAC_2910

//MAC_434 replaced by MAC_2911

//MAC_433 replaced by MAC_2911

//MAC_432 replaced by MAC_2910

//MAC_443 replaced by MAC_2911

//MAC_442 replaced by MAC_2911

//MAC_441 replaced by MAC_2910

//MAC_440 replaced by MAC_2911

//MAC_439 replaced by MAC_2911

//MAC_438 replaced by MAC_2910

//MAC_449 replaced by MAC_2911

//MAC_448 replaced by MAC_2911

//MAC_447 replaced by MAC_2910

//MAC_446 replaced by MAC_2911

//MAC_445 replaced by MAC_2911

//MAC_444 replaced by MAC_2910

//MAC_455 replaced by MAC_2911

//MAC_454 replaced by MAC_2911

//MAC_453 replaced by MAC_2910

//MAC_452 replaced by MAC_2911

//MAC_451 replaced by MAC_2911

//MAC_450 replaced by MAC_2910

//MAC_461 replaced by MAC_2911

//MAC_460 replaced by MAC_2911

//MAC_459 replaced by MAC_2910

//MAC_458 replaced by MAC_2911

//MAC_457 replaced by MAC_2911

//MAC_456 replaced by MAC_2910

//MAC_467 replaced by MAC_2911

//MAC_466 replaced by MAC_2911

//MAC_465 replaced by MAC_2910

//MAC_464 replaced by MAC_2911

//MAC_463 replaced by MAC_2911

//MAC_462 replaced by MAC_2910

//MAC_473 replaced by MAC_2911

//MAC_472 replaced by MAC_2911

//MAC_471 replaced by MAC_2910

//MAC_470 replaced by MAC_2911

//MAC_469 replaced by MAC_2911

//MAC_468 replaced by MAC_2910

//MAC_479 replaced by MAC_2911

//MAC_478 replaced by MAC_2911

//MAC_477 replaced by MAC_2910

//MAC_476 replaced by MAC_2911

//MAC_475 replaced by MAC_2911

//MAC_474 replaced by MAC_2910

//MAC_485 replaced by MAC_2911

//MAC_484 replaced by MAC_2911

//MAC_483 replaced by MAC_2910

//MAC_482 replaced by MAC_2911

//MAC_481 replaced by MAC_2911

//MAC_480 replaced by MAC_2910

//MAC_491 replaced by MAC_2911

//MAC_490 replaced by MAC_2911

//MAC_489 replaced by MAC_2910

//MAC_488 replaced by MAC_2911

//MAC_487 replaced by MAC_2911

//MAC_486 replaced by MAC_2910

//MAC_497 replaced by MAC_2911

//MAC_496 replaced by MAC_2911

//MAC_495 replaced by MAC_2910

//MAC_494 replaced by MAC_2911

//MAC_493 replaced by MAC_2911

//MAC_492 replaced by MAC_2910

//MAC_503 replaced by MAC_2911

//MAC_502 replaced by MAC_2911

//MAC_501 replaced by MAC_2910

//MAC_500 replaced by MAC_2911

//MAC_499 replaced by MAC_2911

//MAC_498 replaced by MAC_2910

//MAC_509 replaced by MAC_2911

//MAC_508 replaced by MAC_2911

//MAC_507 replaced by MAC_2910

//MAC_506 replaced by MAC_2911

//MAC_505 replaced by MAC_2911

//MAC_504 replaced by MAC_2910

//MAC_515 replaced by MAC_2911

//MAC_514 replaced by MAC_2911

//MAC_513 replaced by MAC_2910

//MAC_512 replaced by MAC_2911

//MAC_511 replaced by MAC_2911

//MAC_510 replaced by MAC_2910

//MAC_521 replaced by MAC_2911

//MAC_520 replaced by MAC_2911

//MAC_519 replaced by MAC_2910

//MAC_518 replaced by MAC_2911

//MAC_517 replaced by MAC_2911

//MAC_516 replaced by MAC_2910

//MAC_527 replaced by MAC_2911

//MAC_526 replaced by MAC_2911

//MAC_525 replaced by MAC_2910

//MAC_524 replaced by MAC_2911

//MAC_523 replaced by MAC_2911

//MAC_522 replaced by MAC_2910

//MAC_533 replaced by MAC_2911

//MAC_532 replaced by MAC_2911

//MAC_531 replaced by MAC_2910

//MAC_530 replaced by MAC_2911

//MAC_529 replaced by MAC_2911

//MAC_528 replaced by MAC_2910

//MAC_539 replaced by MAC_2911

//MAC_538 replaced by MAC_2911

//MAC_537 replaced by MAC_2910

//MAC_536 replaced by MAC_2911

//MAC_535 replaced by MAC_2911

//MAC_534 replaced by MAC_2910

//MAC_545 replaced by MAC_2911

//MAC_544 replaced by MAC_2911

//MAC_543 replaced by MAC_2910

//MAC_542 replaced by MAC_2911

//MAC_541 replaced by MAC_2911

//MAC_540 replaced by MAC_2910

//MAC_551 replaced by MAC_2911

//MAC_550 replaced by MAC_2911

//MAC_549 replaced by MAC_2910

//MAC_548 replaced by MAC_2911

//MAC_547 replaced by MAC_2911

//MAC_546 replaced by MAC_2910

//MAC_557 replaced by MAC_2911

//MAC_556 replaced by MAC_2911

//MAC_555 replaced by MAC_2910

//MAC_554 replaced by MAC_2911

//MAC_553 replaced by MAC_2911

//MAC_552 replaced by MAC_2910

//MAC_563 replaced by MAC_2911

//MAC_562 replaced by MAC_2911

//MAC_561 replaced by MAC_2910

//MAC_560 replaced by MAC_2911

//MAC_559 replaced by MAC_2911

//MAC_558 replaced by MAC_2910

//MAC_569 replaced by MAC_2911

//MAC_568 replaced by MAC_2911

//MAC_567 replaced by MAC_2910

//MAC_566 replaced by MAC_2911

//MAC_565 replaced by MAC_2911

//MAC_564 replaced by MAC_2910

//MAC_575 replaced by MAC_2911

//MAC_574 replaced by MAC_2911

//MAC_573 replaced by MAC_2910

//MAC_572 replaced by MAC_2911

//MAC_571 replaced by MAC_2911

//MAC_570 replaced by MAC_2910

//MAC_581 replaced by MAC_2911

//MAC_580 replaced by MAC_2911

//MAC_579 replaced by MAC_2910

//MAC_578 replaced by MAC_2911

//MAC_577 replaced by MAC_2911

//MAC_576 replaced by MAC_2910

//MAC_587 replaced by MAC_2911

//MAC_586 replaced by MAC_2911

//MAC_585 replaced by MAC_2910

//MAC_584 replaced by MAC_2911

//MAC_583 replaced by MAC_2911

//MAC_582 replaced by MAC_2910

//MAC_593 replaced by MAC_2911

//MAC_592 replaced by MAC_2911

//MAC_591 replaced by MAC_2910

//MAC_590 replaced by MAC_2911

//MAC_589 replaced by MAC_2911

//MAC_588 replaced by MAC_2910

//MAC_599 replaced by MAC_2911

//MAC_598 replaced by MAC_2911

//MAC_597 replaced by MAC_2910

//MAC_596 replaced by MAC_2911

//MAC_595 replaced by MAC_2911

//MAC_594 replaced by MAC_2910

//MAC_605 replaced by MAC_2911

//MAC_604 replaced by MAC_2911

//MAC_603 replaced by MAC_2910

//MAC_602 replaced by MAC_2911

//MAC_601 replaced by MAC_2911

//MAC_600 replaced by MAC_2910

//MAC_611 replaced by MAC_2911

//MAC_610 replaced by MAC_2911

//MAC_609 replaced by MAC_2910

//MAC_608 replaced by MAC_2911

//MAC_607 replaced by MAC_2911

//MAC_606 replaced by MAC_2910

//MAC_617 replaced by MAC_2911

//MAC_616 replaced by MAC_2911

//MAC_615 replaced by MAC_2910

//MAC_614 replaced by MAC_2911

//MAC_613 replaced by MAC_2911

//MAC_612 replaced by MAC_2910

//MAC_623 replaced by MAC_2911

//MAC_622 replaced by MAC_2911

//MAC_621 replaced by MAC_2910

//MAC_620 replaced by MAC_2911

//MAC_619 replaced by MAC_2911

//MAC_618 replaced by MAC_2910

//MAC_629 replaced by MAC_2911

//MAC_628 replaced by MAC_2911

//MAC_627 replaced by MAC_2910

//MAC_626 replaced by MAC_2911

//MAC_625 replaced by MAC_2911

//MAC_624 replaced by MAC_2910

//MAC_635 replaced by MAC_2911

//MAC_634 replaced by MAC_2911

//MAC_633 replaced by MAC_2910

//MAC_632 replaced by MAC_2911

//MAC_631 replaced by MAC_2911

//MAC_630 replaced by MAC_2910

//MAC_641 replaced by MAC_2911

//MAC_640 replaced by MAC_2911

//MAC_639 replaced by MAC_2910

//MAC_638 replaced by MAC_2911

//MAC_637 replaced by MAC_2911

//MAC_636 replaced by MAC_2910

//MAC_647 replaced by MAC_2911

//MAC_646 replaced by MAC_2911

//MAC_645 replaced by MAC_2910

//MAC_644 replaced by MAC_2911

//MAC_643 replaced by MAC_2911

//MAC_642 replaced by MAC_2910

//MAC_653 replaced by MAC_2911

//MAC_652 replaced by MAC_2911

//MAC_651 replaced by MAC_2910

//MAC_650 replaced by MAC_2911

//MAC_649 replaced by MAC_2911

//MAC_648 replaced by MAC_2910

//MAC_659 replaced by MAC_2911

//MAC_658 replaced by MAC_2911

//MAC_657 replaced by MAC_2910

//MAC_656 replaced by MAC_2911

//MAC_655 replaced by MAC_2911

//MAC_654 replaced by MAC_2910

//MAC_665 replaced by MAC_2911

//MAC_664 replaced by MAC_2911

//MAC_663 replaced by MAC_2910

//MAC_662 replaced by MAC_2911

//MAC_661 replaced by MAC_2911

//MAC_660 replaced by MAC_2910

//MAC_671 replaced by MAC_2911

//MAC_670 replaced by MAC_2911

//MAC_669 replaced by MAC_2910

//MAC_668 replaced by MAC_2911

//MAC_667 replaced by MAC_2911

//MAC_666 replaced by MAC_2910

//MAC_677 replaced by MAC_2911

//MAC_676 replaced by MAC_2911

//MAC_675 replaced by MAC_2910

//MAC_674 replaced by MAC_2911

//MAC_673 replaced by MAC_2911

//MAC_672 replaced by MAC_2910

//MAC_683 replaced by MAC_2911

//MAC_682 replaced by MAC_2911

//MAC_681 replaced by MAC_2910

//MAC_680 replaced by MAC_2911

//MAC_679 replaced by MAC_2911

//MAC_678 replaced by MAC_2910

//MAC_689 replaced by MAC_2911

//MAC_688 replaced by MAC_2911

//MAC_687 replaced by MAC_2910

//MAC_686 replaced by MAC_2911

//MAC_685 replaced by MAC_2911

//MAC_684 replaced by MAC_2910

//MAC_695 replaced by MAC_2911

//MAC_694 replaced by MAC_2911

//MAC_693 replaced by MAC_2910

//MAC_692 replaced by MAC_2911

//MAC_691 replaced by MAC_2911

//MAC_690 replaced by MAC_2910

//MAC_701 replaced by MAC_2911

//MAC_700 replaced by MAC_2911

//MAC_699 replaced by MAC_2910

//MAC_698 replaced by MAC_2911

//MAC_697 replaced by MAC_2911

//MAC_696 replaced by MAC_2910

//MAC_707 replaced by MAC_2911

//MAC_706 replaced by MAC_2911

//MAC_705 replaced by MAC_2910

//MAC_704 replaced by MAC_2911

//MAC_703 replaced by MAC_2911

//MAC_702 replaced by MAC_2910

//MAC_713 replaced by MAC_2911

//MAC_712 replaced by MAC_2911

//MAC_711 replaced by MAC_2910

//MAC_710 replaced by MAC_2911

//MAC_709 replaced by MAC_2911

//MAC_708 replaced by MAC_2910

//MAC_719 replaced by MAC_2911

//MAC_718 replaced by MAC_2911

//MAC_717 replaced by MAC_2910

//MAC_716 replaced by MAC_2911

//MAC_715 replaced by MAC_2911

//MAC_714 replaced by MAC_2910

//MAC_725 replaced by MAC_2911

//MAC_724 replaced by MAC_2911

//MAC_723 replaced by MAC_2910

//MAC_722 replaced by MAC_2911

//MAC_721 replaced by MAC_2911

//MAC_720 replaced by MAC_2910

//MAC_731 replaced by MAC_2911

//MAC_730 replaced by MAC_2911

//MAC_729 replaced by MAC_2910

//MAC_728 replaced by MAC_2911

//MAC_727 replaced by MAC_2911

//MAC_726 replaced by MAC_2910

//MAC_737 replaced by MAC_2911

//MAC_736 replaced by MAC_2911

//MAC_735 replaced by MAC_2910

//MAC_734 replaced by MAC_2911

//MAC_733 replaced by MAC_2911

//MAC_732 replaced by MAC_2910

//MAC_743 replaced by MAC_2911

//MAC_742 replaced by MAC_2911

//MAC_741 replaced by MAC_2910

//MAC_740 replaced by MAC_2911

//MAC_739 replaced by MAC_2911

//MAC_738 replaced by MAC_2910

//MAC_749 replaced by MAC_2911

//MAC_748 replaced by MAC_2911

//MAC_747 replaced by MAC_2910

//MAC_746 replaced by MAC_2911

//MAC_745 replaced by MAC_2911

//MAC_744 replaced by MAC_2910

//MAC_755 replaced by MAC_2911

//MAC_754 replaced by MAC_2911

//MAC_753 replaced by MAC_2910

//MAC_752 replaced by MAC_2911

//MAC_751 replaced by MAC_2911

//MAC_750 replaced by MAC_2910

//MAC_761 replaced by MAC_2911

//MAC_760 replaced by MAC_2911

//MAC_759 replaced by MAC_2910

//MAC_758 replaced by MAC_2911

//MAC_757 replaced by MAC_2911

//MAC_756 replaced by MAC_2910

//MAC_767 replaced by MAC_2911

//MAC_766 replaced by MAC_2911

//MAC_765 replaced by MAC_2910

//MAC_764 replaced by MAC_2911

//MAC_763 replaced by MAC_2911

//MAC_762 replaced by MAC_2910

//MAC_773 replaced by MAC_2911

//MAC_772 replaced by MAC_2911

//MAC_771 replaced by MAC_2910

//MAC_770 replaced by MAC_2911

//MAC_769 replaced by MAC_2911

//MAC_768 replaced by MAC_2910

//MAC_779 replaced by MAC_2911

//MAC_778 replaced by MAC_2911

//MAC_777 replaced by MAC_2910

//MAC_776 replaced by MAC_2911

//MAC_775 replaced by MAC_2911

//MAC_774 replaced by MAC_2910

//MAC_785 replaced by MAC_2911

//MAC_784 replaced by MAC_2911

//MAC_783 replaced by MAC_2910

//MAC_782 replaced by MAC_2911

//MAC_781 replaced by MAC_2911

//MAC_780 replaced by MAC_2910

//MAC_791 replaced by MAC_2911

//MAC_790 replaced by MAC_2911

//MAC_789 replaced by MAC_2910

//MAC_788 replaced by MAC_2911

//MAC_787 replaced by MAC_2911

//MAC_786 replaced by MAC_2910

//MAC_797 replaced by MAC_2911

//MAC_796 replaced by MAC_2911

//MAC_795 replaced by MAC_2910

//MAC_794 replaced by MAC_2911

//MAC_793 replaced by MAC_2911

//MAC_792 replaced by MAC_2910

//MAC_803 replaced by MAC_2911

//MAC_802 replaced by MAC_2911

//MAC_801 replaced by MAC_2910

//MAC_800 replaced by MAC_2911

//MAC_799 replaced by MAC_2911

//MAC_798 replaced by MAC_2910

//MAC_809 replaced by MAC_2911

//MAC_808 replaced by MAC_2911

//MAC_807 replaced by MAC_2910

//MAC_806 replaced by MAC_2911

//MAC_805 replaced by MAC_2911

//MAC_804 replaced by MAC_2910

//MAC_815 replaced by MAC_2911

//MAC_814 replaced by MAC_2911

//MAC_813 replaced by MAC_2910

//MAC_812 replaced by MAC_2911

//MAC_811 replaced by MAC_2911

//MAC_810 replaced by MAC_2910

//MAC_821 replaced by MAC_2911

//MAC_820 replaced by MAC_2911

//MAC_819 replaced by MAC_2910

//MAC_818 replaced by MAC_2911

//MAC_817 replaced by MAC_2911

//MAC_816 replaced by MAC_2910

//MAC_827 replaced by MAC_2911

//MAC_826 replaced by MAC_2911

//MAC_825 replaced by MAC_2910

//MAC_824 replaced by MAC_2911

//MAC_823 replaced by MAC_2911

//MAC_822 replaced by MAC_2910

//MAC_833 replaced by MAC_2911

//MAC_832 replaced by MAC_2911

//MAC_831 replaced by MAC_2910

//MAC_830 replaced by MAC_2911

//MAC_829 replaced by MAC_2911

//MAC_828 replaced by MAC_2910

//MAC_839 replaced by MAC_2911

//MAC_838 replaced by MAC_2911

//MAC_837 replaced by MAC_2910

//MAC_836 replaced by MAC_2911

//MAC_835 replaced by MAC_2911

//MAC_834 replaced by MAC_2910

//MAC_845 replaced by MAC_2911

//MAC_844 replaced by MAC_2911

//MAC_843 replaced by MAC_2910

//MAC_842 replaced by MAC_2911

//MAC_841 replaced by MAC_2911

//MAC_840 replaced by MAC_2910

//MAC_851 replaced by MAC_2911

//MAC_850 replaced by MAC_2911

//MAC_849 replaced by MAC_2910

//MAC_848 replaced by MAC_2911

//MAC_847 replaced by MAC_2911

//MAC_846 replaced by MAC_2910

//MAC_857 replaced by MAC_2911

//MAC_856 replaced by MAC_2911

//MAC_855 replaced by MAC_2910

//MAC_854 replaced by MAC_2911

//MAC_853 replaced by MAC_2911

//MAC_852 replaced by MAC_2910

//MAC_863 replaced by MAC_2911

//MAC_862 replaced by MAC_2911

//MAC_861 replaced by MAC_2910

//MAC_860 replaced by MAC_2911

//MAC_859 replaced by MAC_2911

//MAC_858 replaced by MAC_2910

//MAC_869 replaced by MAC_2911

//MAC_868 replaced by MAC_2911

//MAC_867 replaced by MAC_2910

//MAC_866 replaced by MAC_2911

//MAC_865 replaced by MAC_2911

//MAC_864 replaced by MAC_2910

//MAC_875 replaced by MAC_2911

//MAC_874 replaced by MAC_2911

//MAC_873 replaced by MAC_2910

//MAC_872 replaced by MAC_2911

//MAC_871 replaced by MAC_2911

//MAC_870 replaced by MAC_2910

//MAC_881 replaced by MAC_2911

//MAC_880 replaced by MAC_2911

//MAC_879 replaced by MAC_2910

//MAC_878 replaced by MAC_2911

//MAC_877 replaced by MAC_2911

//MAC_876 replaced by MAC_2910

//MAC_887 replaced by MAC_2911

//MAC_886 replaced by MAC_2911

//MAC_885 replaced by MAC_2910

//MAC_884 replaced by MAC_2911

//MAC_883 replaced by MAC_2911

//MAC_882 replaced by MAC_2910

//MAC_893 replaced by MAC_2911

//MAC_892 replaced by MAC_2911

//MAC_891 replaced by MAC_2910

//MAC_890 replaced by MAC_2911

//MAC_889 replaced by MAC_2911

//MAC_888 replaced by MAC_2910

//MAC_899 replaced by MAC_2911

//MAC_898 replaced by MAC_2911

//MAC_897 replaced by MAC_2910

//MAC_896 replaced by MAC_2911

//MAC_895 replaced by MAC_2911

//MAC_894 replaced by MAC_2910

//MAC_905 replaced by MAC_2911

//MAC_904 replaced by MAC_2911

//MAC_903 replaced by MAC_2910

//MAC_902 replaced by MAC_2911

//MAC_901 replaced by MAC_2911

//MAC_900 replaced by MAC_2910

//MAC_911 replaced by MAC_2911

//MAC_910 replaced by MAC_2911

//MAC_909 replaced by MAC_2910

//MAC_908 replaced by MAC_2911

//MAC_907 replaced by MAC_2911

//MAC_906 replaced by MAC_2910

//MAC_917 replaced by MAC_2911

//MAC_916 replaced by MAC_2911

//MAC_915 replaced by MAC_2910

//MAC_914 replaced by MAC_2911

//MAC_913 replaced by MAC_2911

//MAC_912 replaced by MAC_2910

//MAC_923 replaced by MAC_2911

//MAC_922 replaced by MAC_2911

//MAC_921 replaced by MAC_2910

//MAC_920 replaced by MAC_2911

//MAC_919 replaced by MAC_2911

//MAC_918 replaced by MAC_2910

//MAC_929 replaced by MAC_2911

//MAC_928 replaced by MAC_2911

//MAC_927 replaced by MAC_2910

//MAC_926 replaced by MAC_2911

//MAC_925 replaced by MAC_2911

//MAC_924 replaced by MAC_2910

//MAC_935 replaced by MAC_2911

//MAC_934 replaced by MAC_2911

//MAC_933 replaced by MAC_2910

//MAC_932 replaced by MAC_2911

//MAC_931 replaced by MAC_2911

//MAC_930 replaced by MAC_2910

//MAC_941 replaced by MAC_2911

//MAC_940 replaced by MAC_2911

//MAC_939 replaced by MAC_2910

//MAC_938 replaced by MAC_2911

//MAC_937 replaced by MAC_2911

//MAC_936 replaced by MAC_2910

//MAC_947 replaced by MAC_2911

//MAC_946 replaced by MAC_2911

//MAC_945 replaced by MAC_2910

//MAC_944 replaced by MAC_2911

//MAC_943 replaced by MAC_2911

//MAC_942 replaced by MAC_2910

//MAC_953 replaced by MAC_2911

//MAC_952 replaced by MAC_2911

//MAC_951 replaced by MAC_2910

//MAC_950 replaced by MAC_2911

//MAC_949 replaced by MAC_2911

//MAC_948 replaced by MAC_2910

//MAC_959 replaced by MAC_2911

//MAC_958 replaced by MAC_2911

//MAC_957 replaced by MAC_2910

//MAC_956 replaced by MAC_2911

//MAC_955 replaced by MAC_2911

//MAC_954 replaced by MAC_2910

//MAC_965 replaced by MAC_2911

//MAC_964 replaced by MAC_2911

//MAC_963 replaced by MAC_2910

//MAC_962 replaced by MAC_2911

//MAC_961 replaced by MAC_2911

//MAC_960 replaced by MAC_2910

//MAC_971 replaced by MAC_2911

//MAC_970 replaced by MAC_2911

//MAC_969 replaced by MAC_2910

//MAC_968 replaced by MAC_2911

//MAC_967 replaced by MAC_2911

//MAC_966 replaced by MAC_2910

//MAC_977 replaced by MAC_2911

//MAC_976 replaced by MAC_2911

//MAC_975 replaced by MAC_2910

//MAC_974 replaced by MAC_2911

//MAC_973 replaced by MAC_2911

//MAC_972 replaced by MAC_2910

//MAC_983 replaced by MAC_2911

//MAC_982 replaced by MAC_2911

//MAC_981 replaced by MAC_2910

//MAC_980 replaced by MAC_2911

//MAC_979 replaced by MAC_2911

//MAC_978 replaced by MAC_2910

//MAC_989 replaced by MAC_2911

//MAC_988 replaced by MAC_2911

//MAC_987 replaced by MAC_2910

//MAC_986 replaced by MAC_2911

//MAC_985 replaced by MAC_2911

//MAC_984 replaced by MAC_2910

//MAC_995 replaced by MAC_2911

//MAC_994 replaced by MAC_2911

//MAC_993 replaced by MAC_2910

//MAC_992 replaced by MAC_2911

//MAC_991 replaced by MAC_2911

//MAC_990 replaced by MAC_2910

//MAC_1001 replaced by MAC_2911

//MAC_1000 replaced by MAC_2911

//MAC_999 replaced by MAC_2910

//MAC_998 replaced by MAC_2911

//MAC_997 replaced by MAC_2911

//MAC_996 replaced by MAC_2910

//MAC_1007 replaced by MAC_2911

//MAC_1006 replaced by MAC_2911

//MAC_1005 replaced by MAC_2910

//MAC_1004 replaced by MAC_2911

//MAC_1003 replaced by MAC_2911

//MAC_1002 replaced by MAC_2910

//MAC_1013 replaced by MAC_2911

//MAC_1012 replaced by MAC_2911

//MAC_1011 replaced by MAC_2910

//MAC_1010 replaced by MAC_2911

//MAC_1009 replaced by MAC_2911

//MAC_1008 replaced by MAC_2910

//MAC_1019 replaced by MAC_2911

//MAC_1018 replaced by MAC_2911

//MAC_1017 replaced by MAC_2910

//MAC_1016 replaced by MAC_2911

//MAC_1015 replaced by MAC_2911

//MAC_1014 replaced by MAC_2910

//MAC_1025 replaced by MAC_2911

//MAC_1024 replaced by MAC_2911

//MAC_1023 replaced by MAC_2910

//MAC_1022 replaced by MAC_2911

//MAC_1021 replaced by MAC_2911

//MAC_1020 replaced by MAC_2910

//MAC_1031 replaced by MAC_2911

//MAC_1030 replaced by MAC_2911

//MAC_1029 replaced by MAC_2910

//MAC_1028 replaced by MAC_2911

//MAC_1027 replaced by MAC_2911

//MAC_1026 replaced by MAC_2910

//MAC_1037 replaced by MAC_2911

//MAC_1036 replaced by MAC_2911

//MAC_1035 replaced by MAC_2910

//MAC_1034 replaced by MAC_2911

//MAC_1033 replaced by MAC_2911

//MAC_1032 replaced by MAC_2910

//MAC_1043 replaced by MAC_2911

//MAC_1042 replaced by MAC_2911

//MAC_1041 replaced by MAC_2910

//MAC_1040 replaced by MAC_2911

//MAC_1039 replaced by MAC_2911

//MAC_1038 replaced by MAC_2910

//MAC_1049 replaced by MAC_2911

//MAC_1048 replaced by MAC_2911

//MAC_1047 replaced by MAC_2910

//MAC_1046 replaced by MAC_2911

//MAC_1045 replaced by MAC_2911

//MAC_1044 replaced by MAC_2910

//MAC_1055 replaced by MAC_2911

//MAC_1054 replaced by MAC_2911

//MAC_1053 replaced by MAC_2910

//MAC_1052 replaced by MAC_2911

//MAC_1051 replaced by MAC_2911

//MAC_1050 replaced by MAC_2910

//MAC_1061 replaced by MAC_2911

//MAC_1060 replaced by MAC_2911

//MAC_1059 replaced by MAC_2910

//MAC_1058 replaced by MAC_2911

//MAC_1057 replaced by MAC_2911

//MAC_1056 replaced by MAC_2910

//MAC_1067 replaced by MAC_2911

//MAC_1066 replaced by MAC_2911

//MAC_1065 replaced by MAC_2910

//MAC_1064 replaced by MAC_2911

//MAC_1063 replaced by MAC_2911

//MAC_1062 replaced by MAC_2910

//MAC_1073 replaced by MAC_2911

//MAC_1072 replaced by MAC_2911

//MAC_1071 replaced by MAC_2910

//MAC_1070 replaced by MAC_2911

//MAC_1069 replaced by MAC_2911

//MAC_1068 replaced by MAC_2910

//MAC_1079 replaced by MAC_2911

//MAC_1078 replaced by MAC_2911

//MAC_1077 replaced by MAC_2910

//MAC_1076 replaced by MAC_2911

//MAC_1075 replaced by MAC_2911

//MAC_1074 replaced by MAC_2910

//MAC_1085 replaced by MAC_2911

//MAC_1084 replaced by MAC_2911

//MAC_1083 replaced by MAC_2910

//MAC_1082 replaced by MAC_2911

//MAC_1081 replaced by MAC_2911

//MAC_1080 replaced by MAC_2910

//MAC_1091 replaced by MAC_2911

//MAC_1090 replaced by MAC_2911

//MAC_1089 replaced by MAC_2910

//MAC_1088 replaced by MAC_2911

//MAC_1087 replaced by MAC_2911

//MAC_1086 replaced by MAC_2910

//MAC_1097 replaced by MAC_2911

//MAC_1096 replaced by MAC_2911

//MAC_1095 replaced by MAC_2910

//MAC_1094 replaced by MAC_2911

//MAC_1093 replaced by MAC_2911

//MAC_1092 replaced by MAC_2910

//MAC_1103 replaced by MAC_2911

//MAC_1102 replaced by MAC_2911

//MAC_1101 replaced by MAC_2910

//MAC_1100 replaced by MAC_2911

//MAC_1099 replaced by MAC_2911

//MAC_1098 replaced by MAC_2910

//MAC_1109 replaced by MAC_2911

//MAC_1108 replaced by MAC_2911

//MAC_1107 replaced by MAC_2910

//MAC_1106 replaced by MAC_2911

//MAC_1105 replaced by MAC_2911

//MAC_1104 replaced by MAC_2910

//MAC_1115 replaced by MAC_2911

//MAC_1114 replaced by MAC_2911

//MAC_1113 replaced by MAC_2910

//MAC_1112 replaced by MAC_2911

//MAC_1111 replaced by MAC_2911

//MAC_1110 replaced by MAC_2910

//MAC_1121 replaced by MAC_2911

//MAC_1120 replaced by MAC_2911

//MAC_1119 replaced by MAC_2910

//MAC_1118 replaced by MAC_2911

//MAC_1117 replaced by MAC_2911

//MAC_1116 replaced by MAC_2910

//MAC_1127 replaced by MAC_2911

//MAC_1126 replaced by MAC_2911

//MAC_1125 replaced by MAC_2910

//MAC_1124 replaced by MAC_2911

//MAC_1123 replaced by MAC_2911

//MAC_1122 replaced by MAC_2910

//MAC_1133 replaced by MAC_2911

//MAC_1132 replaced by MAC_2911

//MAC_1131 replaced by MAC_2910

//MAC_1130 replaced by MAC_2911

//MAC_1129 replaced by MAC_2911

//MAC_1128 replaced by MAC_2910

//MAC_1139 replaced by MAC_2911

//MAC_1138 replaced by MAC_2911

//MAC_1137 replaced by MAC_2910

//MAC_1136 replaced by MAC_2911

//MAC_1135 replaced by MAC_2911

//MAC_1134 replaced by MAC_2910

//MAC_1145 replaced by MAC_2911

//MAC_1144 replaced by MAC_2911

//MAC_1143 replaced by MAC_2910

//MAC_1142 replaced by MAC_2911

//MAC_1141 replaced by MAC_2911

//MAC_1140 replaced by MAC_2910

//MAC_1151 replaced by MAC_2911

//MAC_1150 replaced by MAC_2911

//MAC_1149 replaced by MAC_2910

//MAC_1148 replaced by MAC_2911

//MAC_1147 replaced by MAC_2911

//MAC_1146 replaced by MAC_2910

//MAC_1157 replaced by MAC_2911

//MAC_1156 replaced by MAC_2911

//MAC_1155 replaced by MAC_2910

//MAC_1154 replaced by MAC_2911

//MAC_1153 replaced by MAC_2911

//MAC_1152 replaced by MAC_2910

//MAC_1163 replaced by MAC_2911

//MAC_1162 replaced by MAC_2911

//MAC_1161 replaced by MAC_2910

//MAC_1160 replaced by MAC_2911

//MAC_1159 replaced by MAC_2911

//MAC_1158 replaced by MAC_2910

//MAC_1169 replaced by MAC_2911

//MAC_1168 replaced by MAC_2911

//MAC_1167 replaced by MAC_2910

//MAC_1166 replaced by MAC_2911

//MAC_1165 replaced by MAC_2911

//MAC_1164 replaced by MAC_2910

//MAC_1175 replaced by MAC_2911

//MAC_1174 replaced by MAC_2911

//MAC_1173 replaced by MAC_2910

//MAC_1172 replaced by MAC_2911

//MAC_1171 replaced by MAC_2911

//MAC_1170 replaced by MAC_2910

//MAC_1181 replaced by MAC_2911

//MAC_1180 replaced by MAC_2911

//MAC_1179 replaced by MAC_2910

//MAC_1178 replaced by MAC_2911

//MAC_1177 replaced by MAC_2911

//MAC_1176 replaced by MAC_2910

//MAC_1187 replaced by MAC_2911

//MAC_1186 replaced by MAC_2911

//MAC_1185 replaced by MAC_2910

//MAC_1184 replaced by MAC_2911

//MAC_1183 replaced by MAC_2911

//MAC_1182 replaced by MAC_2910

//MAC_1193 replaced by MAC_2911

//MAC_1192 replaced by MAC_2911

//MAC_1191 replaced by MAC_2910

//MAC_1190 replaced by MAC_2911

//MAC_1189 replaced by MAC_2911

//MAC_1188 replaced by MAC_2910

//MAC_1199 replaced by MAC_2911

//MAC_1198 replaced by MAC_2911

//MAC_1197 replaced by MAC_2910

//MAC_1196 replaced by MAC_2911

//MAC_1195 replaced by MAC_2911

//MAC_1194 replaced by MAC_2910

//MAC_1205 replaced by MAC_2911

//MAC_1204 replaced by MAC_2911

//MAC_1203 replaced by MAC_2910

//MAC_1202 replaced by MAC_2911

//MAC_1201 replaced by MAC_2911

//MAC_1200 replaced by MAC_2910

//MAC_1211 replaced by MAC_2911

//MAC_1210 replaced by MAC_2911

//MAC_1209 replaced by MAC_2910

//MAC_1208 replaced by MAC_2911

//MAC_1207 replaced by MAC_2911

//MAC_1206 replaced by MAC_2910

//MAC_1217 replaced by MAC_2911

//MAC_1216 replaced by MAC_2911

//MAC_1215 replaced by MAC_2910

//MAC_1214 replaced by MAC_2911

//MAC_1213 replaced by MAC_2911

//MAC_1212 replaced by MAC_2910

//MAC_1223 replaced by MAC_2911

//MAC_1222 replaced by MAC_2911

//MAC_1221 replaced by MAC_2910

//MAC_1220 replaced by MAC_2911

//MAC_1219 replaced by MAC_2911

//MAC_1218 replaced by MAC_2910

//MAC_1229 replaced by MAC_2911

//MAC_1228 replaced by MAC_2911

//MAC_1227 replaced by MAC_2910

//MAC_1226 replaced by MAC_2911

//MAC_1225 replaced by MAC_2911

//MAC_1224 replaced by MAC_2910

//MAC_1235 replaced by MAC_2911

//MAC_1234 replaced by MAC_2911

//MAC_1233 replaced by MAC_2910

//MAC_1232 replaced by MAC_2911

//MAC_1231 replaced by MAC_2911

//MAC_1230 replaced by MAC_2910

//MAC_1241 replaced by MAC_2911

//MAC_1240 replaced by MAC_2911

//MAC_1239 replaced by MAC_2910

//MAC_1238 replaced by MAC_2911

//MAC_1237 replaced by MAC_2911

//MAC_1236 replaced by MAC_2910

//MAC_1247 replaced by MAC_2911

//MAC_1246 replaced by MAC_2911

//MAC_1245 replaced by MAC_2910

//MAC_1244 replaced by MAC_2911

//MAC_1243 replaced by MAC_2911

//MAC_1242 replaced by MAC_2910

//MAC_1253 replaced by MAC_2911

//MAC_1252 replaced by MAC_2911

//MAC_1251 replaced by MAC_2910

//MAC_1250 replaced by MAC_2911

//MAC_1249 replaced by MAC_2911

//MAC_1248 replaced by MAC_2910

//MAC_1259 replaced by MAC_2911

//MAC_1258 replaced by MAC_2911

//MAC_1257 replaced by MAC_2910

//MAC_1256 replaced by MAC_2911

//MAC_1255 replaced by MAC_2911

//MAC_1254 replaced by MAC_2910

//MAC_1265 replaced by MAC_2911

//MAC_1264 replaced by MAC_2911

//MAC_1263 replaced by MAC_2910

//MAC_1262 replaced by MAC_2911

//MAC_1261 replaced by MAC_2911

//MAC_1260 replaced by MAC_2910

//MAC_1271 replaced by MAC_2911

//MAC_1270 replaced by MAC_2911

//MAC_1269 replaced by MAC_2910

//MAC_1268 replaced by MAC_2911

//MAC_1267 replaced by MAC_2911

//MAC_1266 replaced by MAC_2910

//MAC_1277 replaced by MAC_2911

//MAC_1276 replaced by MAC_2911

//MAC_1275 replaced by MAC_2910

//MAC_1274 replaced by MAC_2911

//MAC_1273 replaced by MAC_2911

//MAC_1272 replaced by MAC_2910

//MAC_1283 replaced by MAC_2911

//MAC_1282 replaced by MAC_2911

//MAC_1281 replaced by MAC_2910

//MAC_1280 replaced by MAC_2911

//MAC_1279 replaced by MAC_2911

//MAC_1278 replaced by MAC_2910

//MAC_1289 replaced by MAC_2911

//MAC_1288 replaced by MAC_2911

//MAC_1287 replaced by MAC_2910

//MAC_1286 replaced by MAC_2911

//MAC_1285 replaced by MAC_2911

//MAC_1284 replaced by MAC_2910

//MAC_1295 replaced by MAC_2911

//MAC_1294 replaced by MAC_2911

//MAC_1293 replaced by MAC_2910

//MAC_1292 replaced by MAC_2911

//MAC_1291 replaced by MAC_2911

//MAC_1290 replaced by MAC_2910

//MAC_1301 replaced by MAC_2911

//MAC_1300 replaced by MAC_2911

//MAC_1299 replaced by MAC_2910

//MAC_1298 replaced by MAC_2911

//MAC_1297 replaced by MAC_2911

//MAC_1296 replaced by MAC_2910

//MAC_1307 replaced by MAC_2911

//MAC_1306 replaced by MAC_2911

//MAC_1305 replaced by MAC_2910

//MAC_1304 replaced by MAC_2911

//MAC_1303 replaced by MAC_2911

//MAC_1302 replaced by MAC_2910

//MAC_1313 replaced by MAC_2911

//MAC_1312 replaced by MAC_2911

//MAC_1311 replaced by MAC_2910

//MAC_1310 replaced by MAC_2911

//MAC_1309 replaced by MAC_2911

//MAC_1308 replaced by MAC_2910

//MAC_1319 replaced by MAC_2911

//MAC_1318 replaced by MAC_2911

//MAC_1317 replaced by MAC_2910

//MAC_1316 replaced by MAC_2911

//MAC_1315 replaced by MAC_2911

//MAC_1314 replaced by MAC_2910

//MAC_1325 replaced by MAC_2911

//MAC_1324 replaced by MAC_2911

//MAC_1323 replaced by MAC_2910

//MAC_1322 replaced by MAC_2911

//MAC_1321 replaced by MAC_2911

//MAC_1320 replaced by MAC_2910

//MAC_1331 replaced by MAC_2911

//MAC_1330 replaced by MAC_2911

//MAC_1329 replaced by MAC_2910

//MAC_1328 replaced by MAC_2911

//MAC_1327 replaced by MAC_2911

//MAC_1326 replaced by MAC_2910

//MAC_1337 replaced by MAC_2911

//MAC_1336 replaced by MAC_2911

//MAC_1335 replaced by MAC_2910

//MAC_1334 replaced by MAC_2911

//MAC_1333 replaced by MAC_2911

//MAC_1332 replaced by MAC_2910

//MAC_1343 replaced by MAC_2911

//MAC_1342 replaced by MAC_2911

//MAC_1341 replaced by MAC_2910

//MAC_1340 replaced by MAC_2911

//MAC_1339 replaced by MAC_2911

//MAC_1338 replaced by MAC_2910

//MAC_1349 replaced by MAC_2911

//MAC_1348 replaced by MAC_2911

//MAC_1347 replaced by MAC_2910

//MAC_1346 replaced by MAC_2911

//MAC_1345 replaced by MAC_2911

//MAC_1344 replaced by MAC_2910

//MAC_1355 replaced by MAC_2911

//MAC_1354 replaced by MAC_2911

//MAC_1353 replaced by MAC_2910

//MAC_1352 replaced by MAC_2911

//MAC_1351 replaced by MAC_2911

//MAC_1350 replaced by MAC_2910

//MAC_1361 replaced by MAC_2911

//MAC_1360 replaced by MAC_2911

//MAC_1359 replaced by MAC_2910

//MAC_1358 replaced by MAC_2911

//MAC_1357 replaced by MAC_2911

//MAC_1356 replaced by MAC_2910

//MAC_1367 replaced by MAC_2911

//MAC_1366 replaced by MAC_2911

//MAC_1365 replaced by MAC_2910

//MAC_1364 replaced by MAC_2911

//MAC_1363 replaced by MAC_2911

//MAC_1362 replaced by MAC_2910

//MAC_1373 replaced by MAC_2911

//MAC_1372 replaced by MAC_2911

//MAC_1371 replaced by MAC_2910

//MAC_1370 replaced by MAC_2911

//MAC_1369 replaced by MAC_2911

//MAC_1368 replaced by MAC_2910

//MAC_1379 replaced by MAC_2911

//MAC_1378 replaced by MAC_2911

//MAC_1377 replaced by MAC_2910

//MAC_1376 replaced by MAC_2911

//MAC_1375 replaced by MAC_2911

//MAC_1374 replaced by MAC_2910

//MAC_1385 replaced by MAC_2911

//MAC_1384 replaced by MAC_2911

//MAC_1383 replaced by MAC_2910

//MAC_1382 replaced by MAC_2911

//MAC_1381 replaced by MAC_2911

//MAC_1380 replaced by MAC_2910

//MAC_1391 replaced by MAC_2911

//MAC_1390 replaced by MAC_2911

//MAC_1389 replaced by MAC_2910

//MAC_1388 replaced by MAC_2911

//MAC_1387 replaced by MAC_2911

//MAC_1386 replaced by MAC_2910

//MAC_1397 replaced by MAC_2911

//MAC_1396 replaced by MAC_2911

//MAC_1395 replaced by MAC_2910

//MAC_1394 replaced by MAC_2911

//MAC_1393 replaced by MAC_2911

//MAC_1392 replaced by MAC_2910

//MAC_1403 replaced by MAC_2911

//MAC_1402 replaced by MAC_2911

//MAC_1401 replaced by MAC_2910

//MAC_1400 replaced by MAC_2911

//MAC_1399 replaced by MAC_2911

//MAC_1398 replaced by MAC_2910

//MAC_1409 replaced by MAC_2911

//MAC_1408 replaced by MAC_2911

//MAC_1407 replaced by MAC_2910

//MAC_1406 replaced by MAC_2911

//MAC_1405 replaced by MAC_2911

//MAC_1404 replaced by MAC_2910

//MAC_1415 replaced by MAC_2911

//MAC_1414 replaced by MAC_2911

//MAC_1413 replaced by MAC_2910

//MAC_1412 replaced by MAC_2911

//MAC_1411 replaced by MAC_2911

//MAC_1410 replaced by MAC_2910

//MAC_1421 replaced by MAC_2911

//MAC_1420 replaced by MAC_2911

//MAC_1419 replaced by MAC_2910

//MAC_1418 replaced by MAC_2911

//MAC_1417 replaced by MAC_2911

//MAC_1416 replaced by MAC_2910

//MAC_1427 replaced by MAC_2911

//MAC_1426 replaced by MAC_2911

//MAC_1425 replaced by MAC_2910

//MAC_1424 replaced by MAC_2911

//MAC_1423 replaced by MAC_2911

//MAC_1422 replaced by MAC_2910

//MAC_1433 replaced by MAC_2911

//MAC_1432 replaced by MAC_2911

//MAC_1431 replaced by MAC_2910

//MAC_1430 replaced by MAC_2911

//MAC_1429 replaced by MAC_2911

//MAC_1428 replaced by MAC_2910

//MAC_1439 replaced by MAC_2911

//MAC_1438 replaced by MAC_2911

//MAC_1437 replaced by MAC_2910

//MAC_1436 replaced by MAC_2911

//MAC_1435 replaced by MAC_2911

//MAC_1434 replaced by MAC_2910

//MAC_1445 replaced by MAC_2911

//MAC_1444 replaced by MAC_2911

//MAC_1443 replaced by MAC_2910

//MAC_1442 replaced by MAC_2911

//MAC_1441 replaced by MAC_2911

//MAC_1440 replaced by MAC_2910

//MAC_1451 replaced by MAC_2911

//MAC_1450 replaced by MAC_2911

//MAC_1449 replaced by MAC_2910

//MAC_1448 replaced by MAC_2911

//MAC_1447 replaced by MAC_2911

//MAC_1446 replaced by MAC_2910

//MAC_1457 replaced by MAC_2911

//MAC_1456 replaced by MAC_2911

//MAC_1455 replaced by MAC_2910

//MAC_1454 replaced by MAC_2911

//MAC_1453 replaced by MAC_2911

//MAC_1452 replaced by MAC_2910

//MAC_1463 replaced by MAC_2911

//MAC_1462 replaced by MAC_2911

//MAC_1461 replaced by MAC_2910

//MAC_1460 replaced by MAC_2911

//MAC_1459 replaced by MAC_2911

//MAC_1458 replaced by MAC_2910

//MAC_1469 replaced by MAC_2911

//MAC_1468 replaced by MAC_2911

//MAC_1467 replaced by MAC_2910

//MAC_1466 replaced by MAC_2911

//MAC_1465 replaced by MAC_2911

//MAC_1464 replaced by MAC_2910

//MAC_1475 replaced by MAC_2911

//MAC_1474 replaced by MAC_2911

//MAC_1473 replaced by MAC_2910

//MAC_1472 replaced by MAC_2911

//MAC_1471 replaced by MAC_2911

//MAC_1470 replaced by MAC_2910

//MAC_1481 replaced by MAC_2911

//MAC_1480 replaced by MAC_2911

//MAC_1479 replaced by MAC_2910

//MAC_1478 replaced by MAC_2911

//MAC_1477 replaced by MAC_2911

//MAC_1476 replaced by MAC_2910

//MAC_1487 replaced by MAC_2911

//MAC_1486 replaced by MAC_2911

//MAC_1485 replaced by MAC_2910

//MAC_1484 replaced by MAC_2911

//MAC_1483 replaced by MAC_2911

//MAC_1482 replaced by MAC_2910

//MAC_1493 replaced by MAC_2911

//MAC_1492 replaced by MAC_2911

//MAC_1491 replaced by MAC_2910

//MAC_1490 replaced by MAC_2911

//MAC_1489 replaced by MAC_2911

//MAC_1488 replaced by MAC_2910

//MAC_1499 replaced by MAC_2911

//MAC_1498 replaced by MAC_2911

//MAC_1497 replaced by MAC_2910

//MAC_1496 replaced by MAC_2911

//MAC_1495 replaced by MAC_2911

//MAC_1494 replaced by MAC_2910

//MAC_1505 replaced by MAC_2911

//MAC_1504 replaced by MAC_2911

//MAC_1503 replaced by MAC_2910

//MAC_1502 replaced by MAC_2911

//MAC_1501 replaced by MAC_2911

//MAC_1500 replaced by MAC_2910

//MAC_1511 replaced by MAC_2911

//MAC_1510 replaced by MAC_2911

//MAC_1509 replaced by MAC_2910

//MAC_1508 replaced by MAC_2911

//MAC_1507 replaced by MAC_2911

//MAC_1506 replaced by MAC_2910

//MAC_1517 replaced by MAC_2911

//MAC_1516 replaced by MAC_2911

//MAC_1515 replaced by MAC_2910

//MAC_1514 replaced by MAC_2911

//MAC_1513 replaced by MAC_2911

//MAC_1512 replaced by MAC_2910

//MAC_1523 replaced by MAC_2911

//MAC_1522 replaced by MAC_2911

//MAC_1521 replaced by MAC_2910

//MAC_1520 replaced by MAC_2911

//MAC_1519 replaced by MAC_2911

//MAC_1518 replaced by MAC_2910

//MAC_1529 replaced by MAC_2911

//MAC_1528 replaced by MAC_2911

//MAC_1527 replaced by MAC_2910

//MAC_1526 replaced by MAC_2911

//MAC_1525 replaced by MAC_2911

//MAC_1524 replaced by MAC_2910

//MAC_1535 replaced by MAC_2911

//MAC_1534 replaced by MAC_2911

//MAC_1533 replaced by MAC_2910

//MAC_1532 replaced by MAC_2911

//MAC_1531 replaced by MAC_2911

//MAC_1530 replaced by MAC_2910

//MAC_1541 replaced by MAC_2911

//MAC_1540 replaced by MAC_2911

//MAC_1539 replaced by MAC_2910

//MAC_1538 replaced by MAC_2911

//MAC_1537 replaced by MAC_2911

//MAC_1536 replaced by MAC_2910

//MAC_1547 replaced by MAC_2911

//MAC_1546 replaced by MAC_2911

//MAC_1545 replaced by MAC_2910

//MAC_1544 replaced by MAC_2911

//MAC_1543 replaced by MAC_2911

//MAC_1542 replaced by MAC_2910

//MAC_1553 replaced by MAC_2911

//MAC_1552 replaced by MAC_2911

//MAC_1551 replaced by MAC_2910

//MAC_1550 replaced by MAC_2911

//MAC_1549 replaced by MAC_2911

//MAC_1548 replaced by MAC_2910

//MAC_1559 replaced by MAC_2911

//MAC_1558 replaced by MAC_2911

//MAC_1557 replaced by MAC_2910

//MAC_1556 replaced by MAC_2911

//MAC_1555 replaced by MAC_2911

//MAC_1554 replaced by MAC_2910

//MAC_1565 replaced by MAC_2911

//MAC_1564 replaced by MAC_2911

//MAC_1563 replaced by MAC_2910

//MAC_1562 replaced by MAC_2911

//MAC_1561 replaced by MAC_2911

//MAC_1560 replaced by MAC_2910

//MAC_1571 replaced by MAC_2911

//MAC_1570 replaced by MAC_2911

//MAC_1569 replaced by MAC_2910

//MAC_1568 replaced by MAC_2911

//MAC_1567 replaced by MAC_2911

//MAC_1566 replaced by MAC_2910

//MAC_1577 replaced by MAC_2911

//MAC_1576 replaced by MAC_2911

//MAC_1575 replaced by MAC_2910

//MAC_1574 replaced by MAC_2911

//MAC_1573 replaced by MAC_2911

//MAC_1572 replaced by MAC_2910

//MAC_1583 replaced by MAC_2911

//MAC_1582 replaced by MAC_2911

//MAC_1581 replaced by MAC_2910

//MAC_1580 replaced by MAC_2911

//MAC_1579 replaced by MAC_2911

//MAC_1578 replaced by MAC_2910

//MAC_1589 replaced by MAC_2911

//MAC_1588 replaced by MAC_2911

//MAC_1587 replaced by MAC_2910

//MAC_1586 replaced by MAC_2911

//MAC_1585 replaced by MAC_2911

//MAC_1584 replaced by MAC_2910

//MAC_1595 replaced by MAC_2911

//MAC_1594 replaced by MAC_2911

//MAC_1593 replaced by MAC_2910

//MAC_1592 replaced by MAC_2911

//MAC_1591 replaced by MAC_2911

//MAC_1590 replaced by MAC_2910

//MAC_1601 replaced by MAC_2911

//MAC_1600 replaced by MAC_2911

//MAC_1599 replaced by MAC_2910

//MAC_1598 replaced by MAC_2911

//MAC_1597 replaced by MAC_2911

//MAC_1596 replaced by MAC_2910

//MAC_1607 replaced by MAC_2911

//MAC_1606 replaced by MAC_2911

//MAC_1605 replaced by MAC_2910

//MAC_1604 replaced by MAC_2911

//MAC_1603 replaced by MAC_2911

//MAC_1602 replaced by MAC_2910

//MAC_1613 replaced by MAC_2911

//MAC_1612 replaced by MAC_2911

//MAC_1611 replaced by MAC_2910

//MAC_1610 replaced by MAC_2911

//MAC_1609 replaced by MAC_2911

//MAC_1608 replaced by MAC_2910

//MAC_1619 replaced by MAC_2911

//MAC_1618 replaced by MAC_2911

//MAC_1617 replaced by MAC_2910

//MAC_1616 replaced by MAC_2911

//MAC_1615 replaced by MAC_2911

//MAC_1614 replaced by MAC_2910

//MAC_1625 replaced by MAC_2911

//MAC_1624 replaced by MAC_2911

//MAC_1623 replaced by MAC_2910

//MAC_1622 replaced by MAC_2911

//MAC_1621 replaced by MAC_2911

//MAC_1620 replaced by MAC_2910

//MAC_1631 replaced by MAC_2911

//MAC_1630 replaced by MAC_2911

//MAC_1629 replaced by MAC_2910

//MAC_1628 replaced by MAC_2911

//MAC_1627 replaced by MAC_2911

//MAC_1626 replaced by MAC_2910

//MAC_1637 replaced by MAC_2911

//MAC_1636 replaced by MAC_2911

//MAC_1635 replaced by MAC_2910

//MAC_1634 replaced by MAC_2911

//MAC_1633 replaced by MAC_2911

//MAC_1632 replaced by MAC_2910

//MAC_1643 replaced by MAC_2911

//MAC_1642 replaced by MAC_2911

//MAC_1641 replaced by MAC_2910

//MAC_1640 replaced by MAC_2911

//MAC_1639 replaced by MAC_2911

//MAC_1638 replaced by MAC_2910

//MAC_1649 replaced by MAC_2911

//MAC_1648 replaced by MAC_2911

//MAC_1647 replaced by MAC_2910

//MAC_1646 replaced by MAC_2911

//MAC_1645 replaced by MAC_2911

//MAC_1644 replaced by MAC_2910

//MAC_1655 replaced by MAC_2911

//MAC_1654 replaced by MAC_2911

//MAC_1653 replaced by MAC_2910

//MAC_1652 replaced by MAC_2911

//MAC_1651 replaced by MAC_2911

//MAC_1650 replaced by MAC_2910

//MAC_1661 replaced by MAC_2911

//MAC_1660 replaced by MAC_2911

//MAC_1659 replaced by MAC_2910

//MAC_1658 replaced by MAC_2911

//MAC_1657 replaced by MAC_2911

//MAC_1656 replaced by MAC_2910

//MAC_1667 replaced by MAC_2911

//MAC_1666 replaced by MAC_2911

//MAC_1665 replaced by MAC_2910

//MAC_1664 replaced by MAC_2911

//MAC_1663 replaced by MAC_2911

//MAC_1662 replaced by MAC_2910

//MAC_1673 replaced by MAC_2911

//MAC_1672 replaced by MAC_2911

//MAC_1671 replaced by MAC_2910

//MAC_1670 replaced by MAC_2911

//MAC_1669 replaced by MAC_2911

//MAC_1668 replaced by MAC_2910

//MAC_1679 replaced by MAC_2911

//MAC_1678 replaced by MAC_2911

//MAC_1677 replaced by MAC_2910

//MAC_1676 replaced by MAC_2911

//MAC_1675 replaced by MAC_2911

//MAC_1674 replaced by MAC_2910

//MAC_1685 replaced by MAC_2911

//MAC_1684 replaced by MAC_2911

//MAC_1683 replaced by MAC_2910

//MAC_1682 replaced by MAC_2911

//MAC_1681 replaced by MAC_2911

//MAC_1680 replaced by MAC_2910

//MAC_1691 replaced by MAC_2911

//MAC_1690 replaced by MAC_2911

//MAC_1689 replaced by MAC_2910

//MAC_1688 replaced by MAC_2911

//MAC_1687 replaced by MAC_2911

//MAC_1686 replaced by MAC_2910

//MAC_1697 replaced by MAC_2911

//MAC_1696 replaced by MAC_2911

//MAC_1695 replaced by MAC_2910

//MAC_1694 replaced by MAC_2911

//MAC_1693 replaced by MAC_2911

//MAC_1692 replaced by MAC_2910

//MAC_1703 replaced by MAC_2911

//MAC_1702 replaced by MAC_2911

//MAC_1701 replaced by MAC_2910

//MAC_1700 replaced by MAC_2911

//MAC_1699 replaced by MAC_2911

//MAC_1698 replaced by MAC_2910

//MAC_1709 replaced by MAC_2911

//MAC_1708 replaced by MAC_2911

//MAC_1707 replaced by MAC_2910

//MAC_1706 replaced by MAC_2911

//MAC_1705 replaced by MAC_2911

//MAC_1704 replaced by MAC_2910

//MAC_1715 replaced by MAC_2911

//MAC_1714 replaced by MAC_2911

//MAC_1713 replaced by MAC_2910

//MAC_1712 replaced by MAC_2911

//MAC_1711 replaced by MAC_2911

//MAC_1710 replaced by MAC_2910

//MAC_1721 replaced by MAC_2911

//MAC_1720 replaced by MAC_2911

//MAC_1719 replaced by MAC_2910

//MAC_1718 replaced by MAC_2911

//MAC_1717 replaced by MAC_2911

//MAC_1716 replaced by MAC_2910

//MAC_1727 replaced by MAC_2911

//MAC_1726 replaced by MAC_2911

//MAC_1725 replaced by MAC_2910

//MAC_1724 replaced by MAC_2911

//MAC_1723 replaced by MAC_2911

//MAC_1722 replaced by MAC_2910

//MAC_1733 replaced by MAC_2911

//MAC_1732 replaced by MAC_2911

//MAC_1731 replaced by MAC_2910

//MAC_1730 replaced by MAC_2911

//MAC_1729 replaced by MAC_2911

//MAC_1728 replaced by MAC_2910

//MAC_1739 replaced by MAC_2911

//MAC_1738 replaced by MAC_2911

//MAC_1737 replaced by MAC_2910

//MAC_1736 replaced by MAC_2911

//MAC_1735 replaced by MAC_2911

//MAC_1734 replaced by MAC_2910

//MAC_1745 replaced by MAC_2911

//MAC_1744 replaced by MAC_2911

//MAC_1743 replaced by MAC_2910

//MAC_1742 replaced by MAC_2911

//MAC_1741 replaced by MAC_2911

//MAC_1740 replaced by MAC_2910

//MAC_1751 replaced by MAC_2911

//MAC_1750 replaced by MAC_2911

//MAC_1749 replaced by MAC_2910

//MAC_1748 replaced by MAC_2911

//MAC_1747 replaced by MAC_2911

//MAC_1746 replaced by MAC_2910

//MAC_1757 replaced by MAC_2911

//MAC_1756 replaced by MAC_2911

//MAC_1755 replaced by MAC_2910

//MAC_1754 replaced by MAC_2911

//MAC_1753 replaced by MAC_2911

//MAC_1752 replaced by MAC_2910

//MAC_1763 replaced by MAC_2911

//MAC_1762 replaced by MAC_2911

//MAC_1761 replaced by MAC_2910

//MAC_1760 replaced by MAC_2911

//MAC_1759 replaced by MAC_2911

//MAC_1758 replaced by MAC_2910

//MAC_1769 replaced by MAC_2911

//MAC_1768 replaced by MAC_2911

//MAC_1767 replaced by MAC_2910

//MAC_1766 replaced by MAC_2911

//MAC_1765 replaced by MAC_2911

//MAC_1764 replaced by MAC_2910

//MAC_1775 replaced by MAC_2911

//MAC_1774 replaced by MAC_2911

//MAC_1773 replaced by MAC_2910

//MAC_1772 replaced by MAC_2911

//MAC_1771 replaced by MAC_2911

//MAC_1770 replaced by MAC_2910

//MAC_1781 replaced by MAC_2911

//MAC_1780 replaced by MAC_2911

//MAC_1779 replaced by MAC_2910

//MAC_1778 replaced by MAC_2911

//MAC_1777 replaced by MAC_2911

//MAC_1776 replaced by MAC_2910

//MAC_1787 replaced by MAC_2911

//MAC_1786 replaced by MAC_2911

//MAC_1785 replaced by MAC_2910

//MAC_1784 replaced by MAC_2911

//MAC_1783 replaced by MAC_2911

//MAC_1782 replaced by MAC_2910

//MAC_1793 replaced by MAC_2911

//MAC_1792 replaced by MAC_2911

//MAC_1791 replaced by MAC_2910

//MAC_1790 replaced by MAC_2911

//MAC_1789 replaced by MAC_2911

//MAC_1788 replaced by MAC_2910

//MAC_1799 replaced by MAC_2911

//MAC_1798 replaced by MAC_2911

//MAC_1797 replaced by MAC_2910

//MAC_1796 replaced by MAC_2911

//MAC_1795 replaced by MAC_2911

//MAC_1794 replaced by MAC_2910

//MAC_1805 replaced by MAC_2911

//MAC_1804 replaced by MAC_2911

//MAC_1803 replaced by MAC_2910

//MAC_1802 replaced by MAC_2911

//MAC_1801 replaced by MAC_2911

//MAC_1800 replaced by MAC_2910

//MAC_1811 replaced by MAC_2911

//MAC_1810 replaced by MAC_2911

//MAC_1809 replaced by MAC_2910

//MAC_1808 replaced by MAC_2911

//MAC_1807 replaced by MAC_2911

//MAC_1806 replaced by MAC_2910

//MAC_1817 replaced by MAC_2911

//MAC_1816 replaced by MAC_2911

//MAC_1815 replaced by MAC_2910

//MAC_1814 replaced by MAC_2911

//MAC_1813 replaced by MAC_2911

//MAC_1812 replaced by MAC_2910

//MAC_1823 replaced by MAC_2911

//MAC_1822 replaced by MAC_2911

//MAC_1821 replaced by MAC_2910

//MAC_1820 replaced by MAC_2911

//MAC_1819 replaced by MAC_2911

//MAC_1818 replaced by MAC_2910

//MAC_1829 replaced by MAC_2911

//MAC_1828 replaced by MAC_2911

//MAC_1827 replaced by MAC_2910

//MAC_1826 replaced by MAC_2911

//MAC_1825 replaced by MAC_2911

//MAC_1824 replaced by MAC_2910

//MAC_1835 replaced by MAC_2911

//MAC_1834 replaced by MAC_2911

//MAC_1833 replaced by MAC_2910

//MAC_1832 replaced by MAC_2911

//MAC_1831 replaced by MAC_2911

//MAC_1830 replaced by MAC_2910

//MAC_1841 replaced by MAC_2911

//MAC_1840 replaced by MAC_2911

//MAC_1839 replaced by MAC_2910

//MAC_1838 replaced by MAC_2911

//MAC_1837 replaced by MAC_2911

//MAC_1836 replaced by MAC_2910

//MAC_1847 replaced by MAC_2911

//MAC_1846 replaced by MAC_2911

//MAC_1845 replaced by MAC_2910

//MAC_1844 replaced by MAC_2911

//MAC_1843 replaced by MAC_2911

//MAC_1842 replaced by MAC_2910

//MAC_1853 replaced by MAC_2911

//MAC_1852 replaced by MAC_2911

//MAC_1851 replaced by MAC_2910

//MAC_1850 replaced by MAC_2911

//MAC_1849 replaced by MAC_2911

//MAC_1848 replaced by MAC_2910

//MAC_1859 replaced by MAC_2911

//MAC_1858 replaced by MAC_2911

//MAC_1857 replaced by MAC_2910

//MAC_1856 replaced by MAC_2911

//MAC_1855 replaced by MAC_2911

//MAC_1854 replaced by MAC_2910

//MAC_1865 replaced by MAC_2911

//MAC_1864 replaced by MAC_2911

//MAC_1863 replaced by MAC_2910

//MAC_1862 replaced by MAC_2911

//MAC_1861 replaced by MAC_2911

//MAC_1860 replaced by MAC_2910

//MAC_1871 replaced by MAC_2911

//MAC_1870 replaced by MAC_2911

//MAC_1869 replaced by MAC_2910

//MAC_1868 replaced by MAC_2911

//MAC_1867 replaced by MAC_2911

//MAC_1866 replaced by MAC_2910

//MAC_1877 replaced by MAC_2911

//MAC_1876 replaced by MAC_2911

//MAC_1875 replaced by MAC_2910

//MAC_1874 replaced by MAC_2911

//MAC_1873 replaced by MAC_2911

//MAC_1872 replaced by MAC_2910

//MAC_1883 replaced by MAC_2911

//MAC_1882 replaced by MAC_2911

//MAC_1881 replaced by MAC_2910

//MAC_1880 replaced by MAC_2911

//MAC_1879 replaced by MAC_2911

//MAC_1878 replaced by MAC_2910

//MAC_1889 replaced by MAC_2911

//MAC_1888 replaced by MAC_2911

//MAC_1887 replaced by MAC_2910

//MAC_1886 replaced by MAC_2911

//MAC_1885 replaced by MAC_2911

//MAC_1884 replaced by MAC_2910

//MAC_1895 replaced by MAC_2911

//MAC_1894 replaced by MAC_2911

//MAC_1893 replaced by MAC_2910

//MAC_1892 replaced by MAC_2911

//MAC_1891 replaced by MAC_2911

//MAC_1890 replaced by MAC_2910

//MAC_1901 replaced by MAC_2911

//MAC_1900 replaced by MAC_2911

//MAC_1899 replaced by MAC_2910

//MAC_1898 replaced by MAC_2911

//MAC_1897 replaced by MAC_2911

//MAC_1896 replaced by MAC_2910

//MAC_1907 replaced by MAC_2911

//MAC_1906 replaced by MAC_2911

//MAC_1905 replaced by MAC_2910

//MAC_1904 replaced by MAC_2911

//MAC_1903 replaced by MAC_2911

//MAC_1902 replaced by MAC_2910

//MAC_1913 replaced by MAC_2911

//MAC_1912 replaced by MAC_2911

//MAC_1911 replaced by MAC_2910

//MAC_1910 replaced by MAC_2911

//MAC_1909 replaced by MAC_2911

//MAC_1908 replaced by MAC_2910

//MAC_1919 replaced by MAC_2911

//MAC_1918 replaced by MAC_2911

//MAC_1917 replaced by MAC_2910

//MAC_1916 replaced by MAC_2911

//MAC_1915 replaced by MAC_2911

//MAC_1914 replaced by MAC_2910

//MAC_1925 replaced by MAC_2911

//MAC_1924 replaced by MAC_2911

//MAC_1923 replaced by MAC_2910

//MAC_1922 replaced by MAC_2911

//MAC_1921 replaced by MAC_2911

//MAC_1920 replaced by MAC_2910

//MAC_1931 replaced by MAC_2911

//MAC_1930 replaced by MAC_2911

//MAC_1929 replaced by MAC_2910

//MAC_1928 replaced by MAC_2911

//MAC_1927 replaced by MAC_2911

//MAC_1926 replaced by MAC_2910

//MAC_1937 replaced by MAC_2911

//MAC_1936 replaced by MAC_2911

//MAC_1935 replaced by MAC_2910

//MAC_1934 replaced by MAC_2911

//MAC_1933 replaced by MAC_2911

//MAC_1932 replaced by MAC_2910

//MAC_1943 replaced by MAC_2911

//MAC_1942 replaced by MAC_2911

//MAC_1941 replaced by MAC_2910

//MAC_1940 replaced by MAC_2911

//MAC_1939 replaced by MAC_2911

//MAC_1938 replaced by MAC_2910

//MAC_1949 replaced by MAC_2911

//MAC_1948 replaced by MAC_2911

//MAC_1947 replaced by MAC_2910

//MAC_1946 replaced by MAC_2911

//MAC_1945 replaced by MAC_2911

//MAC_1944 replaced by MAC_2910

//MAC_1955 replaced by MAC_2911

//MAC_1954 replaced by MAC_2911

//MAC_1953 replaced by MAC_2910

//MAC_1952 replaced by MAC_2911

//MAC_1951 replaced by MAC_2911

//MAC_1950 replaced by MAC_2910

//MAC_1961 replaced by MAC_2911

//MAC_1960 replaced by MAC_2911

//MAC_1959 replaced by MAC_2910

//MAC_1958 replaced by MAC_2911

//MAC_1957 replaced by MAC_2911

//MAC_1956 replaced by MAC_2910

//MAC_1967 replaced by MAC_2911

//MAC_1966 replaced by MAC_2911

//MAC_1965 replaced by MAC_2910

//MAC_1964 replaced by MAC_2911

//MAC_1963 replaced by MAC_2911

//MAC_1962 replaced by MAC_2910

//MAC_1973 replaced by MAC_2911

//MAC_1972 replaced by MAC_2911

//MAC_1971 replaced by MAC_2910

//MAC_1970 replaced by MAC_2911

//MAC_1969 replaced by MAC_2911

//MAC_1968 replaced by MAC_2910

//MAC_1979 replaced by MAC_2911

//MAC_1978 replaced by MAC_2911

//MAC_1977 replaced by MAC_2910

//MAC_1976 replaced by MAC_2911

//MAC_1975 replaced by MAC_2911

//MAC_1974 replaced by MAC_2910

//MAC_1985 replaced by MAC_2911

//MAC_1984 replaced by MAC_2911

//MAC_1983 replaced by MAC_2910

//MAC_1982 replaced by MAC_2911

//MAC_1981 replaced by MAC_2911

//MAC_1980 replaced by MAC_2910

//MAC_1991 replaced by MAC_2911

//MAC_1990 replaced by MAC_2911

//MAC_1989 replaced by MAC_2910

//MAC_1988 replaced by MAC_2911

//MAC_1987 replaced by MAC_2911

//MAC_1986 replaced by MAC_2910

//MAC_1997 replaced by MAC_2911

//MAC_1996 replaced by MAC_2911

//MAC_1995 replaced by MAC_2910

//MAC_1994 replaced by MAC_2911

//MAC_1993 replaced by MAC_2911

//MAC_1992 replaced by MAC_2910

//MAC_2003 replaced by MAC_2911

//MAC_2002 replaced by MAC_2911

//MAC_2001 replaced by MAC_2910

//MAC_2000 replaced by MAC_2911

//MAC_1999 replaced by MAC_2911

//MAC_1998 replaced by MAC_2910

//MAC_2009 replaced by MAC_2911

//MAC_2008 replaced by MAC_2911

//MAC_2007 replaced by MAC_2910

//MAC_2006 replaced by MAC_2911

//MAC_2005 replaced by MAC_2911

//MAC_2004 replaced by MAC_2910

//MAC_2015 replaced by MAC_2911

//MAC_2014 replaced by MAC_2911

//MAC_2013 replaced by MAC_2910

//MAC_2012 replaced by MAC_2911

//MAC_2011 replaced by MAC_2911

//MAC_2010 replaced by MAC_2910

//MAC_2021 replaced by MAC_2911

//MAC_2020 replaced by MAC_2911

//MAC_2019 replaced by MAC_2910

//MAC_2018 replaced by MAC_2911

//MAC_2017 replaced by MAC_2911

//MAC_2016 replaced by MAC_2910

//MAC_2027 replaced by MAC_2911

//MAC_2026 replaced by MAC_2911

//MAC_2025 replaced by MAC_2910

//MAC_2024 replaced by MAC_2911

//MAC_2023 replaced by MAC_2911

//MAC_2022 replaced by MAC_2910

//MAC_2033 replaced by MAC_2911

//MAC_2032 replaced by MAC_2911

//MAC_2031 replaced by MAC_2910

//MAC_2030 replaced by MAC_2911

//MAC_2029 replaced by MAC_2911

//MAC_2028 replaced by MAC_2910

//MAC_2039 replaced by MAC_2911

//MAC_2038 replaced by MAC_2911

//MAC_2037 replaced by MAC_2910

//MAC_2036 replaced by MAC_2911

//MAC_2035 replaced by MAC_2911

//MAC_2034 replaced by MAC_2910

//MAC_2045 replaced by MAC_2911

//MAC_2044 replaced by MAC_2911

//MAC_2043 replaced by MAC_2910

//MAC_2042 replaced by MAC_2911

//MAC_2041 replaced by MAC_2911

//MAC_2040 replaced by MAC_2910

//MAC_2051 replaced by MAC_2911

//MAC_2050 replaced by MAC_2911

//MAC_2049 replaced by MAC_2910

//MAC_2048 replaced by MAC_2911

//MAC_2047 replaced by MAC_2911

//MAC_2046 replaced by MAC_2910

//MAC_2057 replaced by MAC_2911

//MAC_2056 replaced by MAC_2911

//MAC_2055 replaced by MAC_2910

//MAC_2054 replaced by MAC_2911

//MAC_2053 replaced by MAC_2911

//MAC_2052 replaced by MAC_2910

//MAC_2063 replaced by MAC_2911

//MAC_2062 replaced by MAC_2911

//MAC_2061 replaced by MAC_2910

//MAC_2060 replaced by MAC_2911

//MAC_2059 replaced by MAC_2911

//MAC_2058 replaced by MAC_2910

//MAC_2069 replaced by MAC_2911

//MAC_2068 replaced by MAC_2911

//MAC_2067 replaced by MAC_2910

//MAC_2066 replaced by MAC_2911

//MAC_2065 replaced by MAC_2911

//MAC_2064 replaced by MAC_2910

//MAC_2075 replaced by MAC_2911

//MAC_2074 replaced by MAC_2911

//MAC_2073 replaced by MAC_2910

//MAC_2072 replaced by MAC_2911

//MAC_2071 replaced by MAC_2911

//MAC_2070 replaced by MAC_2910

//MAC_2081 replaced by MAC_2911

//MAC_2080 replaced by MAC_2911

//MAC_2079 replaced by MAC_2910

//MAC_2078 replaced by MAC_2911

//MAC_2077 replaced by MAC_2911

//MAC_2076 replaced by MAC_2910

//MAC_2087 replaced by MAC_2911

//MAC_2086 replaced by MAC_2911

//MAC_2085 replaced by MAC_2910

//MAC_2084 replaced by MAC_2911

//MAC_2083 replaced by MAC_2911

//MAC_2082 replaced by MAC_2910

//MAC_2093 replaced by MAC_2911

//MAC_2092 replaced by MAC_2911

//MAC_2091 replaced by MAC_2910

//MAC_2090 replaced by MAC_2911

//MAC_2089 replaced by MAC_2911

//MAC_2088 replaced by MAC_2910

//MAC_2099 replaced by MAC_2911

//MAC_2098 replaced by MAC_2911

//MAC_2097 replaced by MAC_2910

//MAC_2096 replaced by MAC_2911

//MAC_2095 replaced by MAC_2911

//MAC_2094 replaced by MAC_2910

//MAC_2105 replaced by MAC_2911

//MAC_2104 replaced by MAC_2911

//MAC_2103 replaced by MAC_2910

//MAC_2102 replaced by MAC_2911

//MAC_2101 replaced by MAC_2911

//MAC_2100 replaced by MAC_2910

//MAC_2111 replaced by MAC_2911

//MAC_2110 replaced by MAC_2911

//MAC_2109 replaced by MAC_2910

//MAC_2108 replaced by MAC_2911

//MAC_2107 replaced by MAC_2911

//MAC_2106 replaced by MAC_2910

//MAC_2117 replaced by MAC_2911

//MAC_2116 replaced by MAC_2911

//MAC_2115 replaced by MAC_2910

//MAC_2114 replaced by MAC_2911

//MAC_2113 replaced by MAC_2911

//MAC_2112 replaced by MAC_2910

//MAC_2123 replaced by MAC_2911

//MAC_2122 replaced by MAC_2911

//MAC_2121 replaced by MAC_2910

//MAC_2120 replaced by MAC_2911

//MAC_2119 replaced by MAC_2911

//MAC_2118 replaced by MAC_2910

//MAC_2129 replaced by MAC_2911

//MAC_2128 replaced by MAC_2911

//MAC_2127 replaced by MAC_2910

//MAC_2126 replaced by MAC_2911

//MAC_2125 replaced by MAC_2911

//MAC_2124 replaced by MAC_2910

//MAC_2135 replaced by MAC_2911

//MAC_2134 replaced by MAC_2911

//MAC_2133 replaced by MAC_2910

//MAC_2132 replaced by MAC_2911

//MAC_2131 replaced by MAC_2911

//MAC_2130 replaced by MAC_2910

//MAC_2141 replaced by MAC_2911

//MAC_2140 replaced by MAC_2911

//MAC_2139 replaced by MAC_2910

//MAC_2138 replaced by MAC_2911

//MAC_2137 replaced by MAC_2911

//MAC_2136 replaced by MAC_2910

//MAC_2147 replaced by MAC_2911

//MAC_2146 replaced by MAC_2911

//MAC_2145 replaced by MAC_2910

//MAC_2144 replaced by MAC_2911

//MAC_2143 replaced by MAC_2911

//MAC_2142 replaced by MAC_2910

//MAC_2153 replaced by MAC_2911

//MAC_2152 replaced by MAC_2911

//MAC_2151 replaced by MAC_2910

//MAC_2150 replaced by MAC_2911

//MAC_2149 replaced by MAC_2911

//MAC_2148 replaced by MAC_2910

//MAC_2159 replaced by MAC_2911

//MAC_2158 replaced by MAC_2911

//MAC_2157 replaced by MAC_2910

//MAC_2156 replaced by MAC_2911

//MAC_2155 replaced by MAC_2911

//MAC_2154 replaced by MAC_2910

//MAC_2165 replaced by MAC_2911

//MAC_2164 replaced by MAC_2911

//MAC_2163 replaced by MAC_2910

//MAC_2162 replaced by MAC_2911

//MAC_2161 replaced by MAC_2911

//MAC_2160 replaced by MAC_2910

//MAC_2171 replaced by MAC_2911

//MAC_2170 replaced by MAC_2911

//MAC_2169 replaced by MAC_2910

//MAC_2168 replaced by MAC_2911

//MAC_2167 replaced by MAC_2911

//MAC_2166 replaced by MAC_2910

//MAC_2177 replaced by MAC_2911

//MAC_2176 replaced by MAC_2911

//MAC_2175 replaced by MAC_2910

//MAC_2174 replaced by MAC_2911

//MAC_2173 replaced by MAC_2911

//MAC_2172 replaced by MAC_2910

//MAC_2183 replaced by MAC_2911

//MAC_2182 replaced by MAC_2911

//MAC_2181 replaced by MAC_2910

//MAC_2180 replaced by MAC_2911

//MAC_2179 replaced by MAC_2911

//MAC_2178 replaced by MAC_2910

//MAC_2189 replaced by MAC_2911

//MAC_2188 replaced by MAC_2911

//MAC_2187 replaced by MAC_2910

//MAC_2186 replaced by MAC_2911

//MAC_2185 replaced by MAC_2911

//MAC_2184 replaced by MAC_2910

//MAC_2195 replaced by MAC_2911

//MAC_2194 replaced by MAC_2911

//MAC_2193 replaced by MAC_2910

//MAC_2192 replaced by MAC_2911

//MAC_2191 replaced by MAC_2911

//MAC_2190 replaced by MAC_2910

//MAC_2201 replaced by MAC_2911

//MAC_2200 replaced by MAC_2911

//MAC_2199 replaced by MAC_2910

//MAC_2198 replaced by MAC_2911

//MAC_2197 replaced by MAC_2911

//MAC_2196 replaced by MAC_2910

//MAC_2207 replaced by MAC_2911

//MAC_2206 replaced by MAC_2911

//MAC_2205 replaced by MAC_2910

//MAC_2204 replaced by MAC_2911

//MAC_2203 replaced by MAC_2911

//MAC_2202 replaced by MAC_2910

//MAC_2213 replaced by MAC_2911

//MAC_2212 replaced by MAC_2911

//MAC_2211 replaced by MAC_2910

//MAC_2210 replaced by MAC_2911

//MAC_2209 replaced by MAC_2911

//MAC_2208 replaced by MAC_2910

//MAC_2219 replaced by MAC_2911

//MAC_2218 replaced by MAC_2911

//MAC_2217 replaced by MAC_2910

//MAC_2216 replaced by MAC_2911

//MAC_2215 replaced by MAC_2911

//MAC_2214 replaced by MAC_2910

//MAC_2225 replaced by MAC_2911

//MAC_2224 replaced by MAC_2911

//MAC_2223 replaced by MAC_2910

//MAC_2222 replaced by MAC_2911

//MAC_2221 replaced by MAC_2911

//MAC_2220 replaced by MAC_2910

//MAC_2231 replaced by MAC_2911

//MAC_2230 replaced by MAC_2911

//MAC_2229 replaced by MAC_2910

//MAC_2228 replaced by MAC_2911

//MAC_2227 replaced by MAC_2911

//MAC_2226 replaced by MAC_2910

//MAC_2237 replaced by MAC_2911

//MAC_2236 replaced by MAC_2911

//MAC_2235 replaced by MAC_2910

//MAC_2234 replaced by MAC_2911

//MAC_2233 replaced by MAC_2911

//MAC_2232 replaced by MAC_2910

//MAC_2243 replaced by MAC_2911

//MAC_2242 replaced by MAC_2911

//MAC_2241 replaced by MAC_2910

//MAC_2240 replaced by MAC_2911

//MAC_2239 replaced by MAC_2911

//MAC_2238 replaced by MAC_2910

//MAC_2249 replaced by MAC_2911

//MAC_2248 replaced by MAC_2911

//MAC_2247 replaced by MAC_2910

//MAC_2246 replaced by MAC_2911

//MAC_2245 replaced by MAC_2911

//MAC_2244 replaced by MAC_2910

//MAC_2255 replaced by MAC_2911

//MAC_2254 replaced by MAC_2911

//MAC_2253 replaced by MAC_2910

//MAC_2252 replaced by MAC_2911

//MAC_2251 replaced by MAC_2911

//MAC_2250 replaced by MAC_2910

//MAC_2261 replaced by MAC_2911

//MAC_2260 replaced by MAC_2911

//MAC_2259 replaced by MAC_2910

//MAC_2258 replaced by MAC_2911

//MAC_2257 replaced by MAC_2911

//MAC_2256 replaced by MAC_2910

//MAC_2267 replaced by MAC_2911

//MAC_2266 replaced by MAC_2911

//MAC_2265 replaced by MAC_2910

//MAC_2264 replaced by MAC_2911

//MAC_2263 replaced by MAC_2911

//MAC_2262 replaced by MAC_2910

//MAC_2273 replaced by MAC_2911

//MAC_2272 replaced by MAC_2911

//MAC_2271 replaced by MAC_2910

//MAC_2270 replaced by MAC_2911

//MAC_2269 replaced by MAC_2911

//MAC_2268 replaced by MAC_2910

//MAC_2279 replaced by MAC_2911

//MAC_2278 replaced by MAC_2911

//MAC_2277 replaced by MAC_2910

//MAC_2276 replaced by MAC_2911

//MAC_2275 replaced by MAC_2911

//MAC_2274 replaced by MAC_2910

//MAC_2285 replaced by MAC_2911

//MAC_2284 replaced by MAC_2911

//MAC_2283 replaced by MAC_2910

//MAC_2282 replaced by MAC_2911

//MAC_2281 replaced by MAC_2911

//MAC_2280 replaced by MAC_2910

//MAC_2291 replaced by MAC_2911

//MAC_2290 replaced by MAC_2911

//MAC_2289 replaced by MAC_2910

//MAC_2288 replaced by MAC_2911

//MAC_2287 replaced by MAC_2911

//MAC_2286 replaced by MAC_2910

//MAC_2297 replaced by MAC_2911

//MAC_2296 replaced by MAC_2911

//MAC_2295 replaced by MAC_2910

//MAC_2294 replaced by MAC_2911

//MAC_2293 replaced by MAC_2911

//MAC_2292 replaced by MAC_2910

//MAC_2303 replaced by MAC_2911

//MAC_2302 replaced by MAC_2911

//MAC_2301 replaced by MAC_2910

//MAC_2300 replaced by MAC_2911

//MAC_2299 replaced by MAC_2911

//MAC_2298 replaced by MAC_2910

//MAC_2309 replaced by MAC_2911

//MAC_2308 replaced by MAC_2911

//MAC_2307 replaced by MAC_2910

//MAC_2306 replaced by MAC_2911

//MAC_2305 replaced by MAC_2911

//MAC_2304 replaced by MAC_2910

//MAC_2315 replaced by MAC_2911

//MAC_2314 replaced by MAC_2911

//MAC_2313 replaced by MAC_2910

//MAC_2312 replaced by MAC_2911

//MAC_2311 replaced by MAC_2911

//MAC_2310 replaced by MAC_2910

//MAC_2321 replaced by MAC_2911

//MAC_2320 replaced by MAC_2911

//MAC_2319 replaced by MAC_2910

//MAC_2318 replaced by MAC_2911

//MAC_2317 replaced by MAC_2911

//MAC_2316 replaced by MAC_2910

//MAC_2327 replaced by MAC_2911

//MAC_2326 replaced by MAC_2911

//MAC_2325 replaced by MAC_2910

//MAC_2324 replaced by MAC_2911

//MAC_2323 replaced by MAC_2911

//MAC_2322 replaced by MAC_2910

//MAC_2333 replaced by MAC_2911

//MAC_2332 replaced by MAC_2911

//MAC_2331 replaced by MAC_2910

//MAC_2330 replaced by MAC_2911

//MAC_2329 replaced by MAC_2911

//MAC_2328 replaced by MAC_2910

//MAC_2339 replaced by MAC_2911

//MAC_2338 replaced by MAC_2911

//MAC_2337 replaced by MAC_2910

//MAC_2336 replaced by MAC_2911

//MAC_2335 replaced by MAC_2911

//MAC_2334 replaced by MAC_2910

//MAC_2345 replaced by MAC_2911

//MAC_2344 replaced by MAC_2911

//MAC_2343 replaced by MAC_2910

//MAC_2342 replaced by MAC_2911

//MAC_2341 replaced by MAC_2911

//MAC_2340 replaced by MAC_2910

//MAC_2351 replaced by MAC_2911

//MAC_2350 replaced by MAC_2911

//MAC_2349 replaced by MAC_2910

//MAC_2348 replaced by MAC_2911

//MAC_2347 replaced by MAC_2911

//MAC_2346 replaced by MAC_2910

//MAC_2357 replaced by MAC_2911

//MAC_2356 replaced by MAC_2911

//MAC_2355 replaced by MAC_2910

//MAC_2354 replaced by MAC_2911

//MAC_2353 replaced by MAC_2911

//MAC_2352 replaced by MAC_2910

//MAC_2363 replaced by MAC_2911

//MAC_2362 replaced by MAC_2911

//MAC_2361 replaced by MAC_2910

//MAC_2360 replaced by MAC_2911

//MAC_2359 replaced by MAC_2911

//MAC_2358 replaced by MAC_2910

//MAC_2369 replaced by MAC_2911

//MAC_2368 replaced by MAC_2911

//MAC_2367 replaced by MAC_2910

//MAC_2366 replaced by MAC_2911

//MAC_2365 replaced by MAC_2911

//MAC_2364 replaced by MAC_2910

//MAC_2375 replaced by MAC_2911

//MAC_2374 replaced by MAC_2911

//MAC_2373 replaced by MAC_2910

//MAC_2372 replaced by MAC_2911

//MAC_2371 replaced by MAC_2911

//MAC_2370 replaced by MAC_2910

//MAC_2381 replaced by MAC_2911

//MAC_2380 replaced by MAC_2911

//MAC_2379 replaced by MAC_2910

//MAC_2378 replaced by MAC_2911

//MAC_2377 replaced by MAC_2911

//MAC_2376 replaced by MAC_2910

//MAC_2387 replaced by MAC_2911

//MAC_2386 replaced by MAC_2911

//MAC_2385 replaced by MAC_2910

//MAC_2384 replaced by MAC_2911

//MAC_2383 replaced by MAC_2911

//MAC_2382 replaced by MAC_2910

//MAC_2393 replaced by MAC_2911

//MAC_2392 replaced by MAC_2911

//MAC_2391 replaced by MAC_2910

//MAC_2390 replaced by MAC_2911

//MAC_2389 replaced by MAC_2911

//MAC_2388 replaced by MAC_2910

//MAC_2399 replaced by MAC_2911

//MAC_2398 replaced by MAC_2911

//MAC_2397 replaced by MAC_2910

//MAC_2396 replaced by MAC_2911

//MAC_2395 replaced by MAC_2911

//MAC_2394 replaced by MAC_2910

//MAC_2405 replaced by MAC_2911

//MAC_2404 replaced by MAC_2911

//MAC_2403 replaced by MAC_2910

//MAC_2402 replaced by MAC_2911

//MAC_2401 replaced by MAC_2911

//MAC_2400 replaced by MAC_2910

//MAC_2411 replaced by MAC_2911

//MAC_2410 replaced by MAC_2911

//MAC_2409 replaced by MAC_2910

//MAC_2408 replaced by MAC_2911

//MAC_2407 replaced by MAC_2911

//MAC_2406 replaced by MAC_2910

//MAC_2417 replaced by MAC_2911

//MAC_2416 replaced by MAC_2911

//MAC_2415 replaced by MAC_2910

//MAC_2414 replaced by MAC_2911

//MAC_2413 replaced by MAC_2911

//MAC_2412 replaced by MAC_2910

//MAC_2423 replaced by MAC_2911

//MAC_2422 replaced by MAC_2911

//MAC_2421 replaced by MAC_2910

//MAC_2420 replaced by MAC_2911

//MAC_2419 replaced by MAC_2911

//MAC_2418 replaced by MAC_2910

//MAC_2429 replaced by MAC_2911

//MAC_2428 replaced by MAC_2911

//MAC_2427 replaced by MAC_2910

//MAC_2426 replaced by MAC_2911

//MAC_2425 replaced by MAC_2911

//MAC_2424 replaced by MAC_2910

//MAC_2435 replaced by MAC_2911

//MAC_2434 replaced by MAC_2911

//MAC_2433 replaced by MAC_2910

//MAC_2432 replaced by MAC_2911

//MAC_2431 replaced by MAC_2911

//MAC_2430 replaced by MAC_2910

//MAC_2441 replaced by MAC_2911

//MAC_2440 replaced by MAC_2911

//MAC_2439 replaced by MAC_2910

//MAC_2438 replaced by MAC_2911

//MAC_2437 replaced by MAC_2911

//MAC_2436 replaced by MAC_2910

//MAC_2447 replaced by MAC_2911

//MAC_2446 replaced by MAC_2911

//MAC_2445 replaced by MAC_2910

//MAC_2444 replaced by MAC_2911

//MAC_2443 replaced by MAC_2911

//MAC_2442 replaced by MAC_2910

//MAC_2453 replaced by MAC_2911

//MAC_2452 replaced by MAC_2911

//MAC_2451 replaced by MAC_2910

//MAC_2450 replaced by MAC_2911

//MAC_2449 replaced by MAC_2911

//MAC_2448 replaced by MAC_2910

//MAC_2459 replaced by MAC_2911

//MAC_2458 replaced by MAC_2911

//MAC_2457 replaced by MAC_2910

//MAC_2456 replaced by MAC_2911

//MAC_2455 replaced by MAC_2911

//MAC_2454 replaced by MAC_2910

//MAC_2465 replaced by MAC_2911

//MAC_2464 replaced by MAC_2911

//MAC_2463 replaced by MAC_2910

//MAC_2462 replaced by MAC_2911

//MAC_2461 replaced by MAC_2911

//MAC_2460 replaced by MAC_2910

//MAC_2471 replaced by MAC_2911

//MAC_2470 replaced by MAC_2911

//MAC_2469 replaced by MAC_2910

//MAC_2468 replaced by MAC_2911

//MAC_2467 replaced by MAC_2911

//MAC_2466 replaced by MAC_2910

//MAC_2477 replaced by MAC_2911

//MAC_2476 replaced by MAC_2911

//MAC_2475 replaced by MAC_2910

//MAC_2474 replaced by MAC_2911

//MAC_2473 replaced by MAC_2911

//MAC_2472 replaced by MAC_2910

//MAC_2483 replaced by MAC_2911

//MAC_2482 replaced by MAC_2911

//MAC_2481 replaced by MAC_2910

//MAC_2480 replaced by MAC_2911

//MAC_2479 replaced by MAC_2911

//MAC_2478 replaced by MAC_2910

//MAC_2489 replaced by MAC_2911

//MAC_2488 replaced by MAC_2911

//MAC_2487 replaced by MAC_2910

//MAC_2486 replaced by MAC_2911

//MAC_2485 replaced by MAC_2911

//MAC_2484 replaced by MAC_2910

//MAC_2495 replaced by MAC_2911

//MAC_2494 replaced by MAC_2911

//MAC_2493 replaced by MAC_2910

//MAC_2492 replaced by MAC_2911

//MAC_2491 replaced by MAC_2911

//MAC_2490 replaced by MAC_2910

//MAC_2501 replaced by MAC_2911

//MAC_2500 replaced by MAC_2911

//MAC_2499 replaced by MAC_2910

//MAC_2498 replaced by MAC_2911

//MAC_2497 replaced by MAC_2911

//MAC_2496 replaced by MAC_2910

//MAC_2507 replaced by MAC_2911

//MAC_2506 replaced by MAC_2911

//MAC_2505 replaced by MAC_2910

//MAC_2504 replaced by MAC_2911

//MAC_2503 replaced by MAC_2911

//MAC_2502 replaced by MAC_2910

//MAC_2513 replaced by MAC_2911

//MAC_2512 replaced by MAC_2911

//MAC_2511 replaced by MAC_2910

//MAC_2510 replaced by MAC_2911

//MAC_2509 replaced by MAC_2911

//MAC_2508 replaced by MAC_2910

//MAC_2519 replaced by MAC_2911

//MAC_2518 replaced by MAC_2911

//MAC_2517 replaced by MAC_2910

//MAC_2516 replaced by MAC_2911

//MAC_2515 replaced by MAC_2911

//MAC_2514 replaced by MAC_2910

//MAC_2525 replaced by MAC_2911

//MAC_2524 replaced by MAC_2911

//MAC_2523 replaced by MAC_2910

//MAC_2522 replaced by MAC_2911

//MAC_2521 replaced by MAC_2911

//MAC_2520 replaced by MAC_2910

//MAC_2531 replaced by MAC_2911

//MAC_2530 replaced by MAC_2911

//MAC_2529 replaced by MAC_2910

//MAC_2528 replaced by MAC_2911

//MAC_2527 replaced by MAC_2911

//MAC_2526 replaced by MAC_2910

//MAC_2537 replaced by MAC_2911

//MAC_2536 replaced by MAC_2911

//MAC_2535 replaced by MAC_2910

//MAC_2534 replaced by MAC_2911

//MAC_2533 replaced by MAC_2911

//MAC_2532 replaced by MAC_2910

//MAC_2543 replaced by MAC_2911

//MAC_2542 replaced by MAC_2911

//MAC_2541 replaced by MAC_2910

//MAC_2540 replaced by MAC_2911

//MAC_2539 replaced by MAC_2911

//MAC_2538 replaced by MAC_2910

//MAC_2549 replaced by MAC_2911

//MAC_2548 replaced by MAC_2911

//MAC_2547 replaced by MAC_2910

//MAC_2546 replaced by MAC_2911

//MAC_2545 replaced by MAC_2911

//MAC_2544 replaced by MAC_2910

//MAC_2555 replaced by MAC_2911

//MAC_2554 replaced by MAC_2911

//MAC_2553 replaced by MAC_2910

//MAC_2552 replaced by MAC_2911

//MAC_2551 replaced by MAC_2911

//MAC_2550 replaced by MAC_2910

//MAC_2561 replaced by MAC_2911

//MAC_2560 replaced by MAC_2911

//MAC_2559 replaced by MAC_2910

//MAC_2558 replaced by MAC_2911

//MAC_2557 replaced by MAC_2911

//MAC_2556 replaced by MAC_2910

//MAC_2567 replaced by MAC_2911

//MAC_2566 replaced by MAC_2911

//MAC_2565 replaced by MAC_2910

//MAC_2564 replaced by MAC_2911

//MAC_2563 replaced by MAC_2911

//MAC_2562 replaced by MAC_2910

//MAC_2573 replaced by MAC_2911

//MAC_2572 replaced by MAC_2911

//MAC_2571 replaced by MAC_2910

//MAC_2570 replaced by MAC_2911

//MAC_2569 replaced by MAC_2911

//MAC_2568 replaced by MAC_2910

//MAC_2579 replaced by MAC_2911

//MAC_2578 replaced by MAC_2911

//MAC_2577 replaced by MAC_2910

//MAC_2576 replaced by MAC_2911

//MAC_2575 replaced by MAC_2911

//MAC_2574 replaced by MAC_2910

//MAC_2585 replaced by MAC_2911

//MAC_2584 replaced by MAC_2911

//MAC_2583 replaced by MAC_2910

//MAC_2582 replaced by MAC_2911

//MAC_2581 replaced by MAC_2911

//MAC_2580 replaced by MAC_2910

//MAC_2591 replaced by MAC_2911

//MAC_2590 replaced by MAC_2911

//MAC_2589 replaced by MAC_2910

//MAC_2588 replaced by MAC_2911

//MAC_2587 replaced by MAC_2911

//MAC_2586 replaced by MAC_2910

//MAC_2597 replaced by MAC_2911

//MAC_2596 replaced by MAC_2911

//MAC_2595 replaced by MAC_2910

//MAC_2594 replaced by MAC_2911

//MAC_2593 replaced by MAC_2911

//MAC_2592 replaced by MAC_2910

//MAC_2603 replaced by MAC_2911

//MAC_2602 replaced by MAC_2911

//MAC_2601 replaced by MAC_2910

//MAC_2600 replaced by MAC_2911

//MAC_2599 replaced by MAC_2911

//MAC_2598 replaced by MAC_2910

//MAC_2609 replaced by MAC_2911

//MAC_2608 replaced by MAC_2911

//MAC_2607 replaced by MAC_2910

//MAC_2606 replaced by MAC_2911

//MAC_2605 replaced by MAC_2911

//MAC_2604 replaced by MAC_2910

//MAC_2615 replaced by MAC_2911

//MAC_2614 replaced by MAC_2911

//MAC_2613 replaced by MAC_2910

//MAC_2612 replaced by MAC_2911

//MAC_2611 replaced by MAC_2911

//MAC_2610 replaced by MAC_2910

//MAC_2621 replaced by MAC_2911

//MAC_2620 replaced by MAC_2911

//MAC_2619 replaced by MAC_2910

//MAC_2618 replaced by MAC_2911

//MAC_2617 replaced by MAC_2911

//MAC_2616 replaced by MAC_2910

//MAC_2627 replaced by MAC_2911

//MAC_2626 replaced by MAC_2911

//MAC_2625 replaced by MAC_2910

//MAC_2624 replaced by MAC_2911

//MAC_2623 replaced by MAC_2911

//MAC_2622 replaced by MAC_2910

//MAC_2633 replaced by MAC_2911

//MAC_2632 replaced by MAC_2911

//MAC_2631 replaced by MAC_2910

//MAC_2630 replaced by MAC_2911

//MAC_2629 replaced by MAC_2911

//MAC_2628 replaced by MAC_2910

//MAC_2639 replaced by MAC_2911

//MAC_2638 replaced by MAC_2911

//MAC_2637 replaced by MAC_2910

//MAC_2636 replaced by MAC_2911

//MAC_2635 replaced by MAC_2911

//MAC_2634 replaced by MAC_2910

//MAC_2645 replaced by MAC_2911

//MAC_2644 replaced by MAC_2911

//MAC_2643 replaced by MAC_2910

//MAC_2642 replaced by MAC_2911

//MAC_2641 replaced by MAC_2911

//MAC_2640 replaced by MAC_2910

//MAC_2651 replaced by MAC_2911

//MAC_2650 replaced by MAC_2911

//MAC_2649 replaced by MAC_2910

//MAC_2648 replaced by MAC_2911

//MAC_2647 replaced by MAC_2911

//MAC_2646 replaced by MAC_2910

//MAC_2657 replaced by MAC_2911

//MAC_2656 replaced by MAC_2911

//MAC_2655 replaced by MAC_2910

//MAC_2654 replaced by MAC_2911

//MAC_2653 replaced by MAC_2911

//MAC_2652 replaced by MAC_2910

//MAC_2663 replaced by MAC_2911

//MAC_2662 replaced by MAC_2911

//MAC_2661 replaced by MAC_2910

//MAC_2660 replaced by MAC_2911

//MAC_2659 replaced by MAC_2911

//MAC_2658 replaced by MAC_2910

//MAC_2669 replaced by MAC_2911

//MAC_2668 replaced by MAC_2911

//MAC_2667 replaced by MAC_2910

//MAC_2666 replaced by MAC_2911

//MAC_2665 replaced by MAC_2911

//MAC_2664 replaced by MAC_2910

//MAC_2675 replaced by MAC_2911

//MAC_2674 replaced by MAC_2911

//MAC_2673 replaced by MAC_2910

//MAC_2672 replaced by MAC_2911

//MAC_2671 replaced by MAC_2911

//MAC_2670 replaced by MAC_2910

//MAC_2681 replaced by MAC_2911

//MAC_2680 replaced by MAC_2911

//MAC_2679 replaced by MAC_2910

//MAC_2678 replaced by MAC_2911

//MAC_2677 replaced by MAC_2911

//MAC_2676 replaced by MAC_2910

//MAC_2687 replaced by MAC_2911

//MAC_2686 replaced by MAC_2911

//MAC_2685 replaced by MAC_2910

//MAC_2684 replaced by MAC_2911

//MAC_2683 replaced by MAC_2911

//MAC_2682 replaced by MAC_2910

//MAC_2693 replaced by MAC_2911

//MAC_2692 replaced by MAC_2911

//MAC_2691 replaced by MAC_2910

//MAC_2690 replaced by MAC_2911

//MAC_2689 replaced by MAC_2911

//MAC_2688 replaced by MAC_2910

//MAC_2699 replaced by MAC_2911

//MAC_2698 replaced by MAC_2911

//MAC_2697 replaced by MAC_2910

//MAC_2696 replaced by MAC_2911

//MAC_2695 replaced by MAC_2911

//MAC_2694 replaced by MAC_2910

//MAC_2705 replaced by MAC_2911

//MAC_2704 replaced by MAC_2911

//MAC_2703 replaced by MAC_2910

//MAC_2702 replaced by MAC_2911

//MAC_2701 replaced by MAC_2911

//MAC_2700 replaced by MAC_2910

//MAC_2711 replaced by MAC_2911

//MAC_2710 replaced by MAC_2911

//MAC_2709 replaced by MAC_2910

//MAC_2708 replaced by MAC_2911

//MAC_2707 replaced by MAC_2911

//MAC_2706 replaced by MAC_2910

//MAC_2717 replaced by MAC_2911

//MAC_2716 replaced by MAC_2911

//MAC_2715 replaced by MAC_2910

//MAC_2714 replaced by MAC_2911

//MAC_2713 replaced by MAC_2911

//MAC_2712 replaced by MAC_2910

//MAC_2723 replaced by MAC_2911

//MAC_2722 replaced by MAC_2911

//MAC_2721 replaced by MAC_2910

//MAC_2720 replaced by MAC_2911

//MAC_2719 replaced by MAC_2911

//MAC_2718 replaced by MAC_2910

//MAC_2729 replaced by MAC_2911

//MAC_2728 replaced by MAC_2911

//MAC_2727 replaced by MAC_2910

//MAC_2726 replaced by MAC_2911

//MAC_2725 replaced by MAC_2911

//MAC_2724 replaced by MAC_2910

//MAC_2735 replaced by MAC_2911

//MAC_2734 replaced by MAC_2911

//MAC_2733 replaced by MAC_2910

//MAC_2732 replaced by MAC_2911

//MAC_2731 replaced by MAC_2911

//MAC_2730 replaced by MAC_2910

//MAC_2741 replaced by MAC_2911

//MAC_2740 replaced by MAC_2911

//MAC_2739 replaced by MAC_2910

//MAC_2738 replaced by MAC_2911

//MAC_2737 replaced by MAC_2911

//MAC_2736 replaced by MAC_2910

//MAC_2747 replaced by MAC_2911

//MAC_2746 replaced by MAC_2911

//MAC_2745 replaced by MAC_2910

//MAC_2744 replaced by MAC_2911

//MAC_2743 replaced by MAC_2911

//MAC_2742 replaced by MAC_2910

//MAC_2753 replaced by MAC_2911

//MAC_2752 replaced by MAC_2911

//MAC_2751 replaced by MAC_2910

//MAC_2750 replaced by MAC_2911

//MAC_2749 replaced by MAC_2911

//MAC_2748 replaced by MAC_2910

//MAC_2759 replaced by MAC_2911

//MAC_2758 replaced by MAC_2911

//MAC_2757 replaced by MAC_2910

//MAC_2756 replaced by MAC_2911

//MAC_2755 replaced by MAC_2911

//MAC_2754 replaced by MAC_2910

//MAC_2765 replaced by MAC_2911

//MAC_2764 replaced by MAC_2911

//MAC_2763 replaced by MAC_2910

//MAC_2762 replaced by MAC_2911

//MAC_2761 replaced by MAC_2911

//MAC_2760 replaced by MAC_2910

//MAC_2771 replaced by MAC_2911

//MAC_2770 replaced by MAC_2911

//MAC_2769 replaced by MAC_2910

//MAC_2768 replaced by MAC_2911

//MAC_2767 replaced by MAC_2911

//MAC_2766 replaced by MAC_2910

//MAC_2777 replaced by MAC_2911

//MAC_2776 replaced by MAC_2911

//MAC_2775 replaced by MAC_2910

//MAC_2774 replaced by MAC_2911

//MAC_2773 replaced by MAC_2911

//MAC_2772 replaced by MAC_2910

//MAC_2783 replaced by MAC_2911

//MAC_2782 replaced by MAC_2911

//MAC_2781 replaced by MAC_2910

//MAC_2780 replaced by MAC_2911

//MAC_2779 replaced by MAC_2911

//MAC_2778 replaced by MAC_2910

//MAC_2789 replaced by MAC_2911

//MAC_2788 replaced by MAC_2911

//MAC_2787 replaced by MAC_2910

//MAC_2786 replaced by MAC_2911

//MAC_2785 replaced by MAC_2911

//MAC_2784 replaced by MAC_2910

//MAC_2795 replaced by MAC_2911

//MAC_2794 replaced by MAC_2911

//MAC_2793 replaced by MAC_2910

//MAC_2792 replaced by MAC_2911

//MAC_2791 replaced by MAC_2911

//MAC_2790 replaced by MAC_2910

//MAC_2801 replaced by MAC_2911

//MAC_2800 replaced by MAC_2911

//MAC_2799 replaced by MAC_2910

//MAC_2798 replaced by MAC_2911

//MAC_2797 replaced by MAC_2911

//MAC_2796 replaced by MAC_2910

//MAC_2807 replaced by MAC_2911

//MAC_2806 replaced by MAC_2911

//MAC_2805 replaced by MAC_2910

//MAC_2804 replaced by MAC_2911

//MAC_2803 replaced by MAC_2911

//MAC_2802 replaced by MAC_2910

//MAC_2813 replaced by MAC_2911

//MAC_2812 replaced by MAC_2911

//MAC_2811 replaced by MAC_2910

//MAC_2810 replaced by MAC_2911

//MAC_2809 replaced by MAC_2911

//MAC_2808 replaced by MAC_2910

//MAC_2819 replaced by MAC_2911

//MAC_2818 replaced by MAC_2911

//MAC_2817 replaced by MAC_2910

//MAC_2816 replaced by MAC_2911

//MAC_2815 replaced by MAC_2911

//MAC_2814 replaced by MAC_2910

//MAC_2825 replaced by MAC_2911

//MAC_2824 replaced by MAC_2911

//MAC_2823 replaced by MAC_2910

//MAC_2822 replaced by MAC_2911

//MAC_2821 replaced by MAC_2911

//MAC_2820 replaced by MAC_2910

//MAC_2831 replaced by MAC_2911

//MAC_2830 replaced by MAC_2911

//MAC_2829 replaced by MAC_2910

//MAC_2828 replaced by MAC_2911

//MAC_2827 replaced by MAC_2911

//MAC_2826 replaced by MAC_2910

//MAC_2837 replaced by MAC_2911

//MAC_2836 replaced by MAC_2911

//MAC_2835 replaced by MAC_2910

//MAC_2834 replaced by MAC_2911

//MAC_2833 replaced by MAC_2911

//MAC_2832 replaced by MAC_2910

//MAC_2843 replaced by MAC_2911

//MAC_2842 replaced by MAC_2911

//MAC_2841 replaced by MAC_2910

//MAC_2840 replaced by MAC_2911

//MAC_2839 replaced by MAC_2911

//MAC_2838 replaced by MAC_2910

//MAC_2849 replaced by MAC_2911

//MAC_2848 replaced by MAC_2911

//MAC_2847 replaced by MAC_2910

//MAC_2846 replaced by MAC_2911

//MAC_2845 replaced by MAC_2911

//MAC_2844 replaced by MAC_2910

//MAC_2855 replaced by MAC_2911

//MAC_2854 replaced by MAC_2911

//MAC_2853 replaced by MAC_2910

//MAC_2852 replaced by MAC_2911

//MAC_2851 replaced by MAC_2911

//MAC_2850 replaced by MAC_2910

//MAC_2861 replaced by MAC_2911

//MAC_2860 replaced by MAC_2911

//MAC_2859 replaced by MAC_2910

//MAC_2858 replaced by MAC_2911

//MAC_2857 replaced by MAC_2911

//MAC_2856 replaced by MAC_2910

//MAC_2867 replaced by MAC_2911

//MAC_2866 replaced by MAC_2911

//MAC_2865 replaced by MAC_2910

//MAC_2864 replaced by MAC_2911

//MAC_2863 replaced by MAC_2911

//MAC_2862 replaced by MAC_2910

//MAC_2873 replaced by MAC_2911

//MAC_2872 replaced by MAC_2911

//MAC_2871 replaced by MAC_2910

//MAC_2870 replaced by MAC_2911

//MAC_2869 replaced by MAC_2911

//MAC_2868 replaced by MAC_2910

//MAC_2879 replaced by MAC_2911

//MAC_2878 replaced by MAC_2911

//MAC_2877 replaced by MAC_2910

//MAC_2876 replaced by MAC_2911

//MAC_2875 replaced by MAC_2911

//MAC_2874 replaced by MAC_2910

//MAC_2885 replaced by MAC_2911

//MAC_2884 replaced by MAC_2911

//MAC_2883 replaced by MAC_2910

//MAC_2882 replaced by MAC_2911

//MAC_2881 replaced by MAC_2911

//MAC_2880 replaced by MAC_2910

//MAC_2891 replaced by MAC_2911

//MAC_2890 replaced by MAC_2911

//MAC_2889 replaced by MAC_2910

//MAC_2888 replaced by MAC_2911

//MAC_2887 replaced by MAC_2911

//MAC_2886 replaced by MAC_2910

//MAC_2897 replaced by MAC_2911

//MAC_2896 replaced by MAC_2911

//MAC_2895 replaced by MAC_2910

//MAC_2894 replaced by MAC_2911

//MAC_2893 replaced by MAC_2911

//MAC_2892 replaced by MAC_2910

//MAC_2903 replaced by MAC_2911

//MAC_2902 replaced by MAC_2911

//MAC_2901 replaced by MAC_2910

//MAC_2900 replaced by MAC_2911

//MAC_2899 replaced by MAC_2911

//MAC_2898 replaced by MAC_2910

//MAC_2909 replaced by MAC_2911

//MAC_2908 replaced by MAC_2911

//MAC_2907 replaced by MAC_2910

//MAC_2906 replaced by MAC_2911

//MAC_2905 replaced by MAC_2911

//MAC_2904 replaced by MAC_2910

//MAC_2915 replaced by MAC_2911

//MAC_2914 replaced by MAC_2911

//MAC_2913 replaced by MAC_2910

//MAC_2912 replaced by MAC_2911

module MAC_2911 (
  input      [25:0]   io_a,
  input      [29:0]   io_acin,
  output     [29:0]   io_acout,
  input      [16:0]   io_b,
  input      [16:0]   io_c,
  input               io_ce,
  input      [47:0]   io_pcin,
  output     [42:0]   io_p,
  output     [47:0]   io_pcout,
  input               clk
);

  wire       [29:0]   DSP_A;
  wire       [17:0]   DSP_B;
  wire       [47:0]   DSP_C;
  wire       [8:0]    DSP_OPMODE;
  wire       [29:0]   DSP_ACOUT;
  wire       [47:0]   DSP_P;
  wire       [47:0]   DSP_PCOUT;
  wire       [26:0]   _zz_A;
  wire       [0:0]    _zz_A_1;
  wire       [0:0]    _zz_B;
  wire       [17:0]   _zz_C;
  wire       [0:0]    _zz_C_1;
  wire       [47:0]   _zz_io_p;

  assign _zz_A = {_zz_A_1,io_a};
  assign _zz_A_1 = 1'b0;
  assign _zz_B = 1'b0;
  assign _zz_C = {_zz_C_1,io_c};
  assign _zz_C_1 = 1'b0;
  assign _zz_io_p = DSP_P;
  DSP48E2 #(
    .A_INPUT("CASCADE"),
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AMULTSEL("A"),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .AUTORESET_PRIORITY("RESET"),
    .B_INPUT ("DIRECT"),
    .BCASCREG(1),
    .BMULTSEL("B"),
    .BREG(1),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'h0),
    .IS_OPMODE_INVERTED(9'h0),
    .IS_RSTA_INVERTED(1'b0),
    .IS_RSTALLCARRYIN_INVERTED(1'b0),
    .IS_RSTALUMODE_INVERTED(1'b0),
    .IS_RSTB_INVERTED(1'b0),
    .IS_RSTC_INVERTED(1'b0),
    .IS_RSTCTRL_INVERTED(1'b0),
    .IS_RSTD_INVERTED(1'b0),
    .IS_RSTINMODE_INVERTED(1'b0),
    .IS_RSTM_INVERTED(1'b0),
    .IS_RSTP_INVERTED(1'b0),
    .MASK(48'h0),
    .MREG(1),
    .OPMODEREG(1),
    .PATTERN(48'h0),
    .PREADDINSEL("A"),
    .PREG(1),
    .RND(48'h0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48"),
    .USE_WIDEXOR("FALSE"),
    .XORSIMD("XOR24_48_96")
  ) DSP (
    .A             (DSP_A[29:0]    ), //i
    .ACIN          (io_acin[29:0]  ), //i
    .ACOUT         (DSP_ACOUT[29:0]), //o
    .B             (DSP_B[17:0]    ), //i
    .C             (DSP_C[47:0]    ), //i
    .CLK           (clk            ), //i
    .OPMODE        (DSP_OPMODE[8:0]), //i
    .P             (DSP_P[47:0]    ), //o
    .PCIN          (io_pcin[47:0]  ), //i
    .PCOUT         (DSP_PCOUT[47:0]), //o
    .ALUMODE       (4'b0000        ), //i
    .BCIN          (18'h0          ), //i
    .CARRYCASCIN   (1'b0           ), //i
    .CARRYIN       (1'b0           ), //i
    .CARRYINSEL    (3'b000         ), //i
    .CEA1          (1'b0           ), //i
    .CEA2          (1'b1           ), //i
    .CEAD          (1'b0           ), //i
    .CEALUMODE     (1'b0           ), //i
    .CEB1          (1'b0           ), //i
    .CEB2          (1'b1           ), //i
    .CEC           (1'b1           ), //i
    .CECARRYIN     (1'b0           ), //i
    .CECTRL        (1'b1           ), //i
    .CED           (1'b0           ), //i
    .CEINMODE      (1'b0           ), //i
    .CEM           (1'b1           ), //i
    .CEP           (1'b1           ), //i
    .D             (27'h0          ), //i
    .INMODE        (5'h0           ), //i
    .MULTSIGNIN    (1'b0           ), //i
    .RSTA          (1'b0           ), //i
    .RSTALLCARRYIN (1'b0           ), //i
    .RSTALUMODE    (1'b0           ), //i
    .RSTB          (1'b0           ), //i
    .RSTC          (1'b0           ), //i
    .RSTCTRL       (1'b0           ), //i
    .RSTD          (1'b0           ), //i
    .RSTINMODE     (1'b0           ), //i
    .RSTM          (1'b0           ), //i
    .RSTP          (1'b0           )  //i
  );
  assign DSP_A = {{3{_zz_A[26]}}, _zz_A};
  assign io_acout = DSP_ACOUT;
  assign DSP_B = {_zz_B,io_b};
  assign DSP_C = {{30{_zz_C[17]}}, _zz_C};
  assign DSP_OPMODE = {{io_ce,io_ce},7'h55};
  assign io_p = _zz_io_p[42:0];
  assign io_pcout = DSP_PCOUT;

endmodule

module MAC_2910 (
  input      [25:0]   io_a,
  input      [29:0]   io_acin,
  output     [29:0]   io_acout,
  input      [16:0]   io_b,
  input      [16:0]   io_c,
  input               io_ce,
  input      [47:0]   io_pcin,
  output     [42:0]   io_p,
  output     [47:0]   io_pcout,
  input               clk
);

  wire       [29:0]   DSP_A;
  wire       [17:0]   DSP_B;
  wire       [47:0]   DSP_C;
  wire       [8:0]    DSP_OPMODE;
  wire       [29:0]   DSP_ACOUT;
  wire       [47:0]   DSP_P;
  wire       [47:0]   DSP_PCOUT;
  wire       [26:0]   _zz_A;
  wire       [0:0]    _zz_A_1;
  wire       [0:0]    _zz_B;
  wire       [17:0]   _zz_C;
  wire       [0:0]    _zz_C_1;
  wire       [47:0]   _zz_io_p;

  assign _zz_A = {_zz_A_1,io_a};
  assign _zz_A_1 = 1'b0;
  assign _zz_B = 1'b0;
  assign _zz_C = {_zz_C_1,io_c};
  assign _zz_C_1 = 1'b0;
  assign _zz_io_p = DSP_P;
  DSP48E2 #(
    .A_INPUT("DIRECT"),
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AMULTSEL("A"),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .AUTORESET_PRIORITY("RESET"),
    .B_INPUT ("DIRECT"),
    .BCASCREG(1),
    .BMULTSEL("B"),
    .BREG(1),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'h0),
    .IS_OPMODE_INVERTED(9'h0),
    .IS_RSTA_INVERTED(1'b0),
    .IS_RSTALLCARRYIN_INVERTED(1'b0),
    .IS_RSTALUMODE_INVERTED(1'b0),
    .IS_RSTB_INVERTED(1'b0),
    .IS_RSTC_INVERTED(1'b0),
    .IS_RSTCTRL_INVERTED(1'b0),
    .IS_RSTD_INVERTED(1'b0),
    .IS_RSTINMODE_INVERTED(1'b0),
    .IS_RSTM_INVERTED(1'b0),
    .IS_RSTP_INVERTED(1'b0),
    .MASK(48'h0),
    .MREG(1),
    .OPMODEREG(1),
    .PATTERN(48'h0),
    .PREADDINSEL("A"),
    .PREG(1),
    .RND(48'h0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48"),
    .USE_WIDEXOR("FALSE"),
    .XORSIMD("XOR24_48_96")
  ) DSP (
    .A             (DSP_A[29:0]    ), //i
    .ACIN          (io_acin[29:0]  ), //i
    .ACOUT         (DSP_ACOUT[29:0]), //o
    .B             (DSP_B[17:0]    ), //i
    .C             (DSP_C[47:0]    ), //i
    .CLK           (clk            ), //i
    .OPMODE        (DSP_OPMODE[8:0]), //i
    .P             (DSP_P[47:0]    ), //o
    .PCIN          (io_pcin[47:0]  ), //i
    .PCOUT         (DSP_PCOUT[47:0]), //o
    .ALUMODE       (4'b0000        ), //i
    .BCIN          (18'h0          ), //i
    .CARRYCASCIN   (1'b0           ), //i
    .CARRYIN       (1'b0           ), //i
    .CARRYINSEL    (3'b000         ), //i
    .CEA1          (1'b0           ), //i
    .CEA2          (1'b1           ), //i
    .CEAD          (1'b0           ), //i
    .CEALUMODE     (1'b0           ), //i
    .CEB1          (1'b0           ), //i
    .CEB2          (1'b1           ), //i
    .CEC           (1'b1           ), //i
    .CECARRYIN     (1'b0           ), //i
    .CECTRL        (1'b1           ), //i
    .CED           (1'b0           ), //i
    .CEINMODE      (1'b0           ), //i
    .CEM           (1'b1           ), //i
    .CEP           (1'b1           ), //i
    .D             (27'h0          ), //i
    .INMODE        (5'h0           ), //i
    .MULTSIGNIN    (1'b0           ), //i
    .RSTA          (1'b0           ), //i
    .RSTALLCARRYIN (1'b0           ), //i
    .RSTALUMODE    (1'b0           ), //i
    .RSTB          (1'b0           ), //i
    .RSTC          (1'b0           ), //i
    .RSTCTRL       (1'b0           ), //i
    .RSTD          (1'b0           ), //i
    .RSTINMODE     (1'b0           ), //i
    .RSTM          (1'b0           ), //i
    .RSTP          (1'b0           )  //i
  );
  assign DSP_A = {{3{_zz_A[26]}}, _zz_A};
  assign io_acout = DSP_ACOUT;
  assign DSP_B = {_zz_B,io_b};
  assign DSP_C = {{30{_zz_C[17]}}, _zz_C};
  assign DSP_OPMODE = {{io_ce,io_ce},7'h05};
  assign io_p = _zz_io_p[42:0];
  assign io_pcout = DSP_PCOUT;

endmodule
